magic
tech sky130A
magscale 1 2
timestamp 1664299617
<< viali >>
rect 2329 15657 2363 15691
rect 5733 15657 5767 15691
rect 4721 15521 4755 15555
rect 1777 15453 1811 15487
rect 2513 15453 2547 15487
rect 2973 15453 3007 15487
rect 3249 15453 3283 15487
rect 4997 15453 5031 15487
rect 5549 15453 5583 15487
rect 8401 15453 8435 15487
rect 8953 15453 8987 15487
rect 3157 15385 3191 15419
rect 8125 15385 8159 15419
rect 1593 15317 1627 15351
rect 3065 15317 3099 15351
rect 6653 15317 6687 15351
rect 9137 15317 9171 15351
rect 6653 15113 6687 15147
rect 2605 15045 2639 15079
rect 8125 15045 8159 15079
rect 1501 14977 1535 15011
rect 1685 14977 1719 15011
rect 2421 14977 2455 15011
rect 3249 14977 3283 15011
rect 3433 14977 3467 15011
rect 4077 14977 4111 15011
rect 8953 14977 8987 15011
rect 5733 14909 5767 14943
rect 8401 14909 8435 14943
rect 2789 14841 2823 14875
rect 5181 14841 5215 14875
rect 1869 14773 1903 14807
rect 3617 14773 3651 14807
rect 4721 14773 4755 14807
rect 9137 14773 9171 14807
rect 4445 14501 4479 14535
rect 2973 14433 3007 14467
rect 5273 14433 5307 14467
rect 3249 14365 3283 14399
rect 3985 14365 4019 14399
rect 4813 14365 4847 14399
rect 7757 14365 7791 14399
rect 8953 14365 8987 14399
rect 4629 14297 4663 14331
rect 7021 14297 7055 14331
rect 9137 14297 9171 14331
rect 1501 14229 1535 14263
rect 3893 14229 3927 14263
rect 8309 14229 8343 14263
rect 9321 14229 9355 14263
rect 5457 14025 5491 14059
rect 5825 13957 5859 13991
rect 1593 13889 1627 13923
rect 3065 13889 3099 13923
rect 4537 13889 4571 13923
rect 4905 13889 4939 13923
rect 5641 13889 5675 13923
rect 7113 13889 7147 13923
rect 8585 13889 8619 13923
rect 2145 13821 2179 13855
rect 6653 13821 6687 13855
rect 8953 13821 8987 13855
rect 2605 13685 2639 13719
rect 9137 13413 9171 13447
rect 4445 13345 4479 13379
rect 7481 13345 7515 13379
rect 3893 13277 3927 13311
rect 5181 13277 5215 13311
rect 5549 13277 5583 13311
rect 7021 13277 7055 13311
rect 8033 13277 8067 13311
rect 8953 13277 8987 13311
rect 1501 13209 1535 13243
rect 2789 13141 2823 13175
rect 8217 13141 8251 13175
rect 8309 12937 8343 12971
rect 1593 12801 1627 12835
rect 2973 12801 3007 12835
rect 4445 12801 4479 12835
rect 5365 12801 5399 12835
rect 6561 12801 6595 12835
rect 9229 12801 9263 12835
rect 2605 12733 2639 12767
rect 5641 12733 5675 12767
rect 6837 12733 6871 12767
rect 2145 12597 2179 12631
rect 4905 12597 4939 12631
rect 9137 12597 9171 12631
rect 2973 12257 3007 12291
rect 3249 12189 3283 12223
rect 3801 12189 3835 12223
rect 3985 12189 4019 12223
rect 4445 12189 4479 12223
rect 4813 12189 4847 12223
rect 6285 12189 6319 12223
rect 7573 12189 7607 12223
rect 8953 12189 8987 12223
rect 9137 12121 9171 12155
rect 1501 12053 1535 12087
rect 3893 12053 3927 12087
rect 6745 12053 6779 12087
rect 8125 12053 8159 12087
rect 9321 12053 9355 12087
rect 8125 11849 8159 11883
rect 9229 11849 9263 11883
rect 5825 11781 5859 11815
rect 8861 11781 8895 11815
rect 8769 11713 8803 11747
rect 9045 11713 9079 11747
rect 3341 11645 3375 11679
rect 3617 11645 3651 11679
rect 4169 11645 4203 11679
rect 6377 11645 6411 11679
rect 6653 11645 6687 11679
rect 1869 11509 1903 11543
rect 2145 11305 2179 11339
rect 2697 11169 2731 11203
rect 4445 11169 4479 11203
rect 1593 11101 1627 11135
rect 8033 11101 8067 11135
rect 8953 11101 8987 11135
rect 3249 11033 3283 11067
rect 5549 11033 5583 11067
rect 7205 11033 7239 11067
rect 7665 11033 7699 11067
rect 7849 11033 7883 11067
rect 4997 10965 5031 10999
rect 9137 10965 9171 10999
rect 4813 10761 4847 10795
rect 5457 10693 5491 10727
rect 1501 10625 1535 10659
rect 2881 10625 2915 10659
rect 4353 10625 4387 10659
rect 5641 10625 5675 10659
rect 6837 10625 6871 10659
rect 8309 10625 8343 10659
rect 9137 10625 9171 10659
rect 2513 10557 2547 10591
rect 8677 10557 8711 10591
rect 9229 10557 9263 10591
rect 5825 10489 5859 10523
rect 2053 10421 2087 10455
rect 6377 10421 6411 10455
rect 2145 10217 2179 10251
rect 8953 10217 8987 10251
rect 9137 10217 9171 10251
rect 1501 10081 1535 10115
rect 2605 10081 2639 10115
rect 4077 10081 4111 10115
rect 8309 10081 8343 10115
rect 3801 10013 3835 10047
rect 6009 10013 6043 10047
rect 6377 10013 6411 10047
rect 7849 10013 7883 10047
rect 9321 9945 9355 9979
rect 3249 9877 3283 9911
rect 5549 9877 5583 9911
rect 8033 9877 8067 9911
rect 9121 9877 9155 9911
rect 7389 9605 7423 9639
rect 9137 9605 9171 9639
rect 3065 9537 3099 9571
rect 3525 9537 3559 9571
rect 5365 9537 5399 9571
rect 6469 9537 6503 9571
rect 1501 9469 1535 9503
rect 2697 9469 2731 9503
rect 3893 9469 3927 9503
rect 5825 9469 5859 9503
rect 6561 9333 6595 9367
rect 6929 9333 6963 9367
rect 4721 9129 4755 9163
rect 1777 8993 1811 9027
rect 4077 8993 4111 9027
rect 7665 8993 7699 9027
rect 1501 8925 1535 8959
rect 5273 8925 5307 8959
rect 7481 8925 7515 8959
rect 9045 8925 9079 8959
rect 3249 8789 3283 8823
rect 6561 8789 6595 8823
rect 9137 8789 9171 8823
rect 5089 8585 5123 8619
rect 5641 8585 5675 8619
rect 6377 8585 6411 8619
rect 9137 8517 9171 8551
rect 1777 8449 1811 8483
rect 2329 8449 2363 8483
rect 3157 8449 3191 8483
rect 4629 8449 4663 8483
rect 5825 8449 5859 8483
rect 6929 8449 6963 8483
rect 2789 8381 2823 8415
rect 8217 8381 8251 8415
rect 9321 8381 9355 8415
rect 3893 7905 3927 7939
rect 1501 7837 1535 7871
rect 7021 7837 7055 7871
rect 8033 7837 8067 7871
rect 8953 7837 8987 7871
rect 3249 7769 3283 7803
rect 5273 7769 5307 7803
rect 9137 7769 9171 7803
rect 4445 7701 4479 7735
rect 7481 7701 7515 7735
rect 9321 7701 9355 7735
rect 5825 7497 5859 7531
rect 9137 7497 9171 7531
rect 1869 7429 1903 7463
rect 3617 7429 3651 7463
rect 4353 7429 4387 7463
rect 8217 7361 8251 7395
rect 9321 7361 9355 7395
rect 4077 7293 4111 7327
rect 6377 7293 6411 7327
rect 6745 7293 6779 7327
rect 8677 7157 8711 7191
rect 1501 6817 1535 6851
rect 1777 6817 1811 6851
rect 3893 6817 3927 6851
rect 5641 6749 5675 6783
rect 6101 6749 6135 6783
rect 6469 6749 6503 6783
rect 7941 6749 7975 6783
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 5365 6681 5399 6715
rect 3249 6613 3283 6647
rect 8401 6613 8435 6647
rect 9321 6613 9355 6647
rect 2329 6409 2363 6443
rect 3249 6409 3283 6443
rect 4997 6273 5031 6307
rect 5825 6273 5859 6307
rect 6929 6273 6963 6307
rect 8401 6273 8435 6307
rect 1777 6205 1811 6239
rect 4721 6205 4755 6239
rect 6561 6205 6595 6239
rect 5641 6069 5675 6103
rect 8861 6069 8895 6103
rect 1777 5865 1811 5899
rect 3065 5865 3099 5899
rect 5549 5865 5583 5899
rect 7021 5865 7055 5899
rect 8309 5865 8343 5899
rect 7573 5797 7607 5831
rect 3801 5729 3835 5763
rect 6377 5729 6411 5763
rect 1593 5661 1627 5695
rect 2513 5661 2547 5695
rect 3249 5661 3283 5695
rect 7757 5661 7791 5695
rect 8401 5661 8435 5695
rect 9229 5661 9263 5695
rect 1409 5593 1443 5627
rect 4077 5593 4111 5627
rect 8953 5593 8987 5627
rect 9137 5593 9171 5627
rect 2329 5525 2363 5559
rect 9045 5525 9079 5559
rect 4077 5321 4111 5355
rect 5825 5321 5859 5355
rect 7297 5321 7331 5355
rect 6377 5253 6411 5287
rect 6561 5253 6595 5287
rect 9229 5253 9263 5287
rect 4169 5185 4203 5219
rect 7205 5185 7239 5219
rect 9137 5185 9171 5219
rect 5181 5117 5215 5151
rect 6745 4981 6779 5015
rect 3617 4777 3651 4811
rect 4721 4777 4755 4811
rect 5273 4777 5307 4811
rect 6745 4777 6779 4811
rect 7389 4777 7423 4811
rect 8401 4777 8435 4811
rect 9229 4777 9263 4811
rect 3525 4573 3559 4607
rect 4537 4573 4571 4607
rect 5181 4573 5215 4607
rect 5365 4573 5399 4607
rect 6193 4573 6227 4607
rect 6837 4573 6871 4607
rect 7297 4573 7331 4607
rect 7481 4573 7515 4607
rect 8585 4573 8619 4607
rect 9045 4573 9079 4607
rect 6009 4437 6043 4471
rect 7021 4233 7055 4267
rect 7573 4233 7607 4267
rect 3709 4097 3743 4131
rect 4813 4097 4847 4131
rect 5641 4097 5675 4131
rect 6101 4097 6135 4131
rect 6285 4097 6319 4131
rect 6837 4097 6871 4131
rect 7021 4097 7055 4131
rect 7665 4097 7699 4131
rect 9045 4097 9079 4131
rect 4077 4029 4111 4063
rect 6193 4029 6227 4063
rect 4905 3961 4939 3995
rect 5457 3893 5491 3927
rect 9229 3893 9263 3927
rect 3617 3689 3651 3723
rect 4353 3689 4387 3723
rect 4997 3689 5031 3723
rect 6009 3689 6043 3723
rect 3525 3485 3559 3519
rect 3709 3485 3743 3519
rect 4169 3485 4203 3519
rect 4905 3485 4939 3519
rect 6101 3485 6135 3519
rect 7021 3485 7055 3519
rect 7205 3485 7239 3519
rect 8217 3485 8251 3519
rect 9045 3485 9079 3519
rect 7205 3349 7239 3383
rect 8309 3349 8343 3383
rect 9229 3349 9263 3383
rect 4813 3145 4847 3179
rect 6193 3145 6227 3179
rect 7205 3145 7239 3179
rect 7849 3145 7883 3179
rect 3985 3077 4019 3111
rect 3617 3009 3651 3043
rect 4721 3009 4755 3043
rect 4905 3009 4939 3043
rect 5365 3009 5399 3043
rect 5549 3009 5583 3043
rect 6009 3009 6043 3043
rect 7021 3009 7055 3043
rect 7665 3009 7699 3043
rect 8493 3009 8527 3043
rect 8677 3009 8711 3043
rect 9137 3009 9171 3043
rect 9321 3009 9355 3043
rect 9229 2873 9263 2907
rect 5457 2805 5491 2839
rect 8585 2805 8619 2839
rect 3617 2601 3651 2635
rect 8585 2601 8619 2635
rect 9137 2601 9171 2635
rect 3525 2397 3559 2431
rect 3709 2397 3743 2431
rect 4905 2397 4939 2431
rect 5917 2397 5951 2431
rect 6101 2397 6135 2431
rect 6561 2397 6595 2431
rect 6745 2397 6779 2431
rect 7205 2397 7239 2431
rect 7389 2397 7423 2431
rect 8677 2397 8711 2431
rect 9321 2397 9355 2431
rect 4721 2261 4755 2295
rect 6009 2261 6043 2295
rect 6745 2261 6779 2295
rect 7297 2261 7331 2295
rect 3709 2057 3743 2091
rect 4353 2057 4387 2091
rect 4997 2057 5031 2091
rect 5641 2057 5675 2091
rect 6745 2057 6779 2091
rect 8677 2057 8711 2091
rect 9229 2057 9263 2091
rect 3525 1921 3559 1955
rect 4169 1921 4203 1955
rect 4813 1921 4847 1955
rect 4997 1921 5031 1955
rect 5457 1921 5491 1955
rect 6101 1921 6135 1955
rect 6285 1921 6319 1955
rect 6745 1921 6779 1955
rect 6929 1921 6963 1955
rect 7389 1921 7423 1955
rect 8493 1921 8527 1955
rect 9321 1921 9355 1955
rect 7481 1785 7515 1819
rect 6193 1717 6227 1751
rect 6653 1513 6687 1547
rect 3617 1309 3651 1343
rect 3709 1309 3743 1343
rect 4169 1309 4203 1343
rect 4813 1309 4847 1343
rect 5917 1309 5951 1343
rect 6101 1309 6135 1343
rect 6745 1309 6779 1343
rect 7389 1309 7423 1343
rect 7297 1241 7331 1275
rect 4353 1173 4387 1207
rect 4905 1173 4939 1207
rect 6009 1173 6043 1207
<< metal1 >>
rect 13630 16668 13636 16720
rect 13688 16708 13694 16720
rect 15286 16708 15292 16720
rect 13688 16680 15292 16708
rect 13688 16668 13694 16680
rect 15286 16668 15292 16680
rect 15344 16668 15350 16720
rect 920 15802 9844 15824
rect 920 15750 2566 15802
rect 2618 15750 2630 15802
rect 2682 15750 2694 15802
rect 2746 15750 2758 15802
rect 2810 15750 2822 15802
rect 2874 15750 7566 15802
rect 7618 15750 7630 15802
rect 7682 15750 7694 15802
rect 7746 15750 7758 15802
rect 7810 15750 7822 15802
rect 7874 15750 9844 15802
rect 920 15728 9844 15750
rect 2317 15691 2375 15697
rect 2317 15657 2329 15691
rect 2363 15688 2375 15691
rect 2406 15688 2412 15700
rect 2363 15660 2412 15688
rect 2363 15657 2375 15660
rect 2317 15651 2375 15657
rect 2406 15648 2412 15660
rect 2464 15648 2470 15700
rect 5718 15688 5724 15700
rect 5679 15660 5724 15688
rect 5718 15648 5724 15660
rect 5776 15648 5782 15700
rect 4706 15552 4712 15564
rect 4667 15524 4712 15552
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 1762 15484 1768 15496
rect 1723 15456 1768 15484
rect 1762 15444 1768 15456
rect 1820 15444 1826 15496
rect 2501 15487 2559 15493
rect 2501 15484 2513 15487
rect 1872 15456 2513 15484
rect 1118 15376 1124 15428
rect 1176 15416 1182 15428
rect 1872 15416 1900 15456
rect 2501 15453 2513 15456
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 3050 15484 3056 15496
rect 3007 15456 3056 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 3237 15487 3295 15493
rect 3237 15453 3249 15487
rect 3283 15484 3295 15487
rect 4062 15484 4068 15496
rect 3283 15456 4068 15484
rect 3283 15453 3295 15456
rect 3237 15447 3295 15453
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15484 5043 15487
rect 5442 15484 5448 15496
rect 5031 15456 5448 15484
rect 5031 15453 5043 15456
rect 4985 15447 5043 15453
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 5537 15487 5595 15493
rect 5537 15453 5549 15487
rect 5583 15484 5595 15487
rect 6178 15484 6184 15496
rect 5583 15456 6184 15484
rect 5583 15453 5595 15456
rect 5537 15447 5595 15453
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 8386 15444 8392 15496
rect 8444 15484 8450 15496
rect 8941 15487 8999 15493
rect 8444 15456 8489 15484
rect 8444 15444 8450 15456
rect 8941 15453 8953 15487
rect 8987 15484 8999 15487
rect 9030 15484 9036 15496
rect 8987 15456 9036 15484
rect 8987 15453 8999 15456
rect 8941 15447 8999 15453
rect 9030 15444 9036 15456
rect 9088 15444 9094 15496
rect 3142 15416 3148 15428
rect 1176 15388 1900 15416
rect 3103 15388 3148 15416
rect 1176 15376 1182 15388
rect 3142 15376 3148 15388
rect 3200 15376 3206 15428
rect 7834 15416 7840 15428
rect 7682 15388 7840 15416
rect 7834 15376 7840 15388
rect 7892 15376 7898 15428
rect 8110 15416 8116 15428
rect 8071 15388 8116 15416
rect 8110 15376 8116 15388
rect 8168 15376 8174 15428
rect 1302 15308 1308 15360
rect 1360 15348 1366 15360
rect 1581 15351 1639 15357
rect 1581 15348 1593 15351
rect 1360 15320 1593 15348
rect 1360 15308 1366 15320
rect 1581 15317 1593 15320
rect 1627 15317 1639 15351
rect 1581 15311 1639 15317
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 3053 15351 3111 15357
rect 3053 15348 3065 15351
rect 2832 15320 3065 15348
rect 2832 15308 2838 15320
rect 3053 15317 3065 15320
rect 3099 15317 3111 15351
rect 3053 15311 3111 15317
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 6641 15351 6699 15357
rect 6641 15348 6653 15351
rect 5408 15320 6653 15348
rect 5408 15308 5414 15320
rect 6641 15317 6653 15320
rect 6687 15317 6699 15351
rect 9122 15348 9128 15360
rect 9083 15320 9128 15348
rect 6641 15311 6699 15317
rect 9122 15308 9128 15320
rect 9180 15308 9186 15360
rect 920 15258 9844 15280
rect 920 15206 3566 15258
rect 3618 15206 3630 15258
rect 3682 15206 3694 15258
rect 3746 15206 3758 15258
rect 3810 15206 3822 15258
rect 3874 15206 8566 15258
rect 8618 15206 8630 15258
rect 8682 15206 8694 15258
rect 8746 15206 8758 15258
rect 8810 15206 8822 15258
rect 8874 15206 9844 15258
rect 13630 15240 13636 15292
rect 13688 15280 13694 15292
rect 16482 15280 16488 15292
rect 13688 15252 16488 15280
rect 13688 15240 13694 15252
rect 16482 15240 16488 15252
rect 16540 15240 16546 15292
rect 920 15184 9844 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1728 15116 2636 15144
rect 1728 15104 1734 15116
rect 934 15036 940 15088
rect 992 15076 998 15088
rect 2608 15085 2636 15116
rect 5534 15104 5540 15156
rect 5592 15144 5598 15156
rect 6641 15147 6699 15153
rect 6641 15144 6653 15147
rect 5592 15116 6653 15144
rect 5592 15104 5598 15116
rect 6641 15113 6653 15116
rect 6687 15113 6699 15147
rect 6641 15107 6699 15113
rect 17908 15104 17914 15156
rect 17966 15144 17972 15156
rect 18782 15144 18788 15156
rect 17966 15116 18788 15144
rect 17966 15104 17972 15116
rect 18782 15104 18788 15116
rect 18840 15104 18846 15156
rect 2593 15079 2651 15085
rect 992 15048 2360 15076
rect 992 15036 998 15048
rect 2332 15020 2360 15048
rect 2593 15045 2605 15079
rect 2639 15076 2651 15079
rect 7834 15076 7840 15088
rect 2639 15048 3464 15076
rect 7682 15048 7840 15076
rect 2639 15045 2651 15048
rect 2593 15039 2651 15045
rect 1489 15011 1547 15017
rect 1489 14977 1501 15011
rect 1535 15008 1547 15011
rect 1578 15008 1584 15020
rect 1535 14980 1584 15008
rect 1535 14977 1547 14980
rect 1489 14971 1547 14977
rect 1578 14968 1584 14980
rect 1636 14968 1642 15020
rect 1670 14968 1676 15020
rect 1728 15008 1734 15020
rect 1728 14980 1773 15008
rect 1728 14968 1734 14980
rect 2314 14968 2320 15020
rect 2372 15008 2378 15020
rect 3436 15017 3464 15048
rect 7834 15036 7840 15048
rect 7892 15036 7898 15088
rect 8113 15079 8171 15085
rect 8113 15045 8125 15079
rect 8159 15076 8171 15079
rect 8202 15076 8208 15088
rect 8159 15048 8208 15076
rect 8159 15045 8171 15048
rect 8113 15039 8171 15045
rect 8202 15036 8208 15048
rect 8260 15036 8266 15088
rect 2409 15011 2467 15017
rect 2409 15008 2421 15011
rect 2372 14980 2421 15008
rect 2372 14968 2378 14980
rect 2409 14977 2421 14980
rect 2455 14977 2467 15011
rect 2409 14971 2467 14977
rect 3237 15011 3295 15017
rect 3237 14977 3249 15011
rect 3283 14977 3295 15011
rect 3237 14971 3295 14977
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 3510 15008 3516 15020
rect 3467 14980 3516 15008
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 1394 14900 1400 14952
rect 1452 14940 1458 14952
rect 3252 14940 3280 14971
rect 3510 14968 3516 14980
rect 3568 14968 3574 15020
rect 4062 15008 4068 15020
rect 4023 14980 4068 15008
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 8938 15008 8944 15020
rect 8899 14980 8944 15008
rect 8938 14968 8944 14980
rect 8996 14968 9002 15020
rect 5718 14940 5724 14952
rect 1452 14912 3280 14940
rect 5679 14912 5724 14940
rect 1452 14900 1458 14912
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 8386 14940 8392 14952
rect 8347 14912 8392 14940
rect 8386 14900 8392 14912
rect 8444 14900 8450 14952
rect 2774 14872 2780 14884
rect 2735 14844 2780 14872
rect 2774 14832 2780 14844
rect 2832 14832 2838 14884
rect 4154 14832 4160 14884
rect 4212 14872 4218 14884
rect 5169 14875 5227 14881
rect 5169 14872 5181 14875
rect 4212 14844 5181 14872
rect 4212 14832 4218 14844
rect 5169 14841 5181 14844
rect 5215 14841 5227 14875
rect 5169 14835 5227 14841
rect 13630 14832 13636 14884
rect 13688 14872 13694 14884
rect 17402 14872 17408 14884
rect 13688 14844 17408 14872
rect 13688 14832 13694 14844
rect 17402 14832 17408 14844
rect 17460 14832 17466 14884
rect 290 14764 296 14816
rect 348 14804 354 14816
rect 1857 14807 1915 14813
rect 1857 14804 1869 14807
rect 348 14776 1869 14804
rect 348 14764 354 14776
rect 1857 14773 1869 14776
rect 1903 14773 1915 14807
rect 1857 14767 1915 14773
rect 3605 14807 3663 14813
rect 3605 14773 3617 14807
rect 3651 14804 3663 14807
rect 4062 14804 4068 14816
rect 3651 14776 4068 14804
rect 3651 14773 3663 14776
rect 3605 14767 3663 14773
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 4522 14764 4528 14816
rect 4580 14804 4586 14816
rect 4709 14807 4767 14813
rect 4709 14804 4721 14807
rect 4580 14776 4721 14804
rect 4580 14764 4586 14776
rect 4709 14773 4721 14776
rect 4755 14773 4767 14807
rect 9122 14804 9128 14816
rect 9083 14776 9128 14804
rect 4709 14767 4767 14773
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 15286 14804 15292 14816
rect 13872 14776 15292 14804
rect 13872 14764 13878 14776
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 920 14714 9844 14736
rect 920 14662 2566 14714
rect 2618 14662 2630 14714
rect 2682 14662 2694 14714
rect 2746 14662 2758 14714
rect 2810 14662 2822 14714
rect 2874 14662 7566 14714
rect 7618 14662 7630 14714
rect 7682 14662 7694 14714
rect 7746 14662 7758 14714
rect 7810 14662 7822 14714
rect 7874 14662 9844 14714
rect 13630 14696 13636 14748
rect 13688 14736 13694 14748
rect 14182 14736 14188 14748
rect 13688 14708 14188 14736
rect 13688 14696 13694 14708
rect 14182 14696 14188 14708
rect 14240 14696 14246 14748
rect 920 14640 9844 14662
rect 13630 14560 13636 14612
rect 13688 14600 13694 14612
rect 14826 14600 14832 14612
rect 13688 14572 14832 14600
rect 13688 14560 13694 14572
rect 14826 14560 14832 14572
rect 14884 14560 14890 14612
rect 3970 14492 3976 14544
rect 4028 14492 4034 14544
rect 4430 14532 4436 14544
rect 4391 14504 4436 14532
rect 4430 14492 4436 14504
rect 4488 14492 4494 14544
rect 2961 14467 3019 14473
rect 2961 14433 2973 14467
rect 3007 14464 3019 14467
rect 3988 14464 4016 14492
rect 5258 14464 5264 14476
rect 3007 14436 4016 14464
rect 5219 14436 5264 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 6886 14436 8340 14464
rect 3234 14356 3240 14408
rect 3292 14396 3298 14408
rect 3970 14396 3976 14408
rect 3292 14368 3337 14396
rect 3931 14368 3976 14396
rect 3292 14356 3298 14368
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 4801 14399 4859 14405
rect 4801 14396 4813 14399
rect 4764 14368 4813 14396
rect 4764 14356 4770 14368
rect 4801 14365 4813 14368
rect 4847 14365 4859 14399
rect 4801 14359 4859 14365
rect 6454 14356 6460 14408
rect 6512 14396 6518 14408
rect 6886 14396 6914 14436
rect 6512 14368 6914 14396
rect 7745 14399 7803 14405
rect 6512 14356 6518 14368
rect 7745 14365 7757 14399
rect 7791 14396 7803 14399
rect 8202 14396 8208 14408
rect 7791 14368 8208 14396
rect 7791 14365 7803 14368
rect 7745 14359 7803 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 8312 14396 8340 14436
rect 8386 14424 8392 14476
rect 8444 14464 8450 14476
rect 15378 14464 15384 14476
rect 8444 14436 15384 14464
rect 8444 14424 8450 14436
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8312 14368 8953 14396
rect 8941 14365 8953 14368
rect 8987 14396 8999 14399
rect 9214 14396 9220 14408
rect 8987 14368 9220 14396
rect 8987 14365 8999 14368
rect 8941 14359 8999 14365
rect 9214 14356 9220 14368
rect 9272 14356 9278 14408
rect 15194 14356 15200 14408
rect 15252 14396 15258 14408
rect 17586 14396 17592 14408
rect 15252 14368 17592 14396
rect 15252 14356 15258 14368
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 2498 14288 2504 14340
rect 2556 14288 2562 14340
rect 3510 14288 3516 14340
rect 3568 14328 3574 14340
rect 4617 14331 4675 14337
rect 4617 14328 4629 14331
rect 3568 14300 4629 14328
rect 3568 14288 3574 14300
rect 4617 14297 4629 14300
rect 4663 14328 4675 14331
rect 5350 14328 5356 14340
rect 4663 14300 5356 14328
rect 4663 14297 4675 14300
rect 4617 14291 4675 14297
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 7009 14331 7067 14337
rect 7009 14297 7021 14331
rect 7055 14328 7067 14331
rect 7374 14328 7380 14340
rect 7055 14300 7380 14328
rect 7055 14297 7067 14300
rect 7009 14291 7067 14297
rect 7374 14288 7380 14300
rect 7432 14288 7438 14340
rect 9125 14331 9183 14337
rect 9125 14297 9137 14331
rect 9171 14328 9183 14331
rect 9398 14328 9404 14340
rect 9171 14300 9404 14328
rect 9171 14297 9183 14300
rect 9125 14291 9183 14297
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 3881 14263 3939 14269
rect 3881 14229 3893 14263
rect 3927 14260 3939 14263
rect 3970 14260 3976 14272
rect 3927 14232 3976 14260
rect 3927 14229 3939 14232
rect 3881 14223 3939 14229
rect 3970 14220 3976 14232
rect 4028 14220 4034 14272
rect 8297 14263 8355 14269
rect 8297 14229 8309 14263
rect 8343 14260 8355 14263
rect 8478 14260 8484 14272
rect 8343 14232 8484 14260
rect 8343 14229 8355 14232
rect 8297 14223 8355 14229
rect 8478 14220 8484 14232
rect 8536 14220 8542 14272
rect 9306 14260 9312 14272
rect 9267 14232 9312 14260
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 920 14170 9844 14192
rect 920 14118 3566 14170
rect 3618 14118 3630 14170
rect 3682 14118 3694 14170
rect 3746 14118 3758 14170
rect 3810 14118 3822 14170
rect 3874 14118 8566 14170
rect 8618 14118 8630 14170
rect 8682 14118 8694 14170
rect 8746 14118 8758 14170
rect 8810 14118 8822 14170
rect 8874 14118 9844 14170
rect 12802 14152 12808 14204
rect 12860 14192 12866 14204
rect 17126 14192 17132 14204
rect 12860 14164 17132 14192
rect 12860 14152 12866 14164
rect 17126 14152 17132 14164
rect 17184 14152 17190 14204
rect 920 14096 9844 14118
rect 5442 14056 5448 14068
rect 5403 14028 5448 14056
rect 5442 14016 5448 14028
rect 5500 14016 5506 14068
rect 9122 14056 9128 14068
rect 7116 14028 9128 14056
rect 4062 13948 4068 14000
rect 4120 13948 4126 14000
rect 5074 13948 5080 14000
rect 5132 13988 5138 14000
rect 5813 13991 5871 13997
rect 5813 13988 5825 13991
rect 5132 13960 5825 13988
rect 5132 13948 5138 13960
rect 5813 13957 5825 13960
rect 5859 13957 5871 13991
rect 5813 13951 5871 13957
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1581 13923 1639 13929
rect 1581 13920 1593 13923
rect 1544 13892 1593 13920
rect 1544 13880 1550 13892
rect 1581 13889 1593 13892
rect 1627 13920 1639 13923
rect 2406 13920 2412 13932
rect 1627 13892 2412 13920
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 3053 13923 3111 13929
rect 3053 13920 3065 13923
rect 2832 13892 3065 13920
rect 2832 13880 2838 13892
rect 3053 13889 3065 13892
rect 3099 13889 3111 13923
rect 4522 13920 4528 13932
rect 4483 13892 4528 13920
rect 3053 13883 3111 13889
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4890 13920 4896 13932
rect 4851 13892 4896 13920
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 5500 13892 5641 13920
rect 5500 13880 5506 13892
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 2179 13824 2728 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 2700 13784 2728 13824
rect 2958 13784 2964 13796
rect 2700 13756 2964 13784
rect 2958 13744 2964 13756
rect 3016 13744 3022 13796
rect 5828 13784 5856 13951
rect 7116 13929 7144 14028
rect 9122 14016 9128 14028
rect 9180 14016 9186 14068
rect 8110 13948 8116 14000
rect 8168 13948 8174 14000
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 8478 13880 8484 13932
rect 8536 13920 8542 13932
rect 8573 13923 8631 13929
rect 8573 13920 8585 13923
rect 8536 13892 8585 13920
rect 8536 13880 8542 13892
rect 8573 13889 8585 13892
rect 8619 13889 8631 13923
rect 8573 13883 8631 13889
rect 6638 13852 6644 13864
rect 6599 13824 6644 13852
rect 6638 13812 6644 13824
rect 6696 13812 6702 13864
rect 8938 13852 8944 13864
rect 8899 13824 8944 13852
rect 8938 13812 8944 13824
rect 8996 13812 9002 13864
rect 5994 13784 6000 13796
rect 5828 13756 6000 13784
rect 5994 13744 6000 13756
rect 6052 13744 6058 13796
rect 1762 13676 1768 13728
rect 1820 13716 1826 13728
rect 2498 13716 2504 13728
rect 1820 13688 2504 13716
rect 1820 13676 1826 13688
rect 2498 13676 2504 13688
rect 2556 13676 2562 13728
rect 2593 13719 2651 13725
rect 2593 13685 2605 13719
rect 2639 13716 2651 13719
rect 3050 13716 3056 13728
rect 2639 13688 3056 13716
rect 2639 13685 2651 13688
rect 2593 13679 2651 13685
rect 3050 13676 3056 13688
rect 3108 13716 3114 13728
rect 8018 13716 8024 13728
rect 3108 13688 8024 13716
rect 3108 13676 3114 13688
rect 8018 13676 8024 13688
rect 8076 13676 8082 13728
rect 920 13626 9844 13648
rect 920 13574 2566 13626
rect 2618 13574 2630 13626
rect 2682 13574 2694 13626
rect 2746 13574 2758 13626
rect 2810 13574 2822 13626
rect 2874 13574 7566 13626
rect 7618 13574 7630 13626
rect 7682 13574 7694 13626
rect 7746 13574 7758 13626
rect 7810 13574 7822 13626
rect 7874 13574 9844 13626
rect 920 13552 9844 13574
rect 13722 13540 13728 13592
rect 13780 13580 13786 13592
rect 16022 13580 16028 13592
rect 13780 13552 16028 13580
rect 13780 13540 13786 13552
rect 16022 13540 16028 13552
rect 16080 13540 16086 13592
rect 17908 13540 17914 13592
rect 17966 13580 17972 13592
rect 18966 13580 18972 13592
rect 17966 13552 18972 13580
rect 17966 13540 17972 13552
rect 18966 13540 18972 13552
rect 19024 13540 19030 13592
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 18322 13512 18328 13524
rect 13872 13484 18328 13512
rect 13872 13472 13878 13484
rect 18322 13472 18328 13484
rect 18380 13472 18386 13524
rect 9125 13447 9183 13453
rect 9125 13413 9137 13447
rect 9171 13444 9183 13447
rect 15746 13444 15752 13456
rect 9171 13416 15752 13444
rect 9171 13413 9183 13416
rect 9125 13407 9183 13413
rect 15746 13404 15752 13416
rect 15804 13404 15810 13456
rect 106 13336 112 13388
rect 164 13376 170 13388
rect 1394 13376 1400 13388
rect 164 13348 1400 13376
rect 164 13336 170 13348
rect 1394 13336 1400 13348
rect 1452 13336 1458 13388
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 5442 13376 5448 13388
rect 4479 13348 5448 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 7469 13379 7527 13385
rect 7469 13345 7481 13379
rect 7515 13376 7527 13379
rect 7515 13348 8064 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 3050 13268 3056 13320
rect 3108 13308 3114 13320
rect 3881 13311 3939 13317
rect 3881 13308 3893 13311
rect 3108 13280 3893 13308
rect 3108 13268 3114 13280
rect 3881 13277 3893 13280
rect 3927 13308 3939 13311
rect 4062 13308 4068 13320
rect 3927 13280 4068 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 5166 13308 5172 13320
rect 5127 13280 5172 13308
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 5534 13308 5540 13320
rect 5495 13280 5540 13308
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 7006 13308 7012 13320
rect 6967 13280 7012 13308
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 8036 13317 8064 13348
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13277 8079 13311
rect 8021 13271 8079 13277
rect 8386 13268 8392 13320
rect 8444 13308 8450 13320
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 8444 13280 8953 13308
rect 8444 13268 8450 13280
rect 8941 13277 8953 13280
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 1394 13200 1400 13252
rect 1452 13240 1458 13252
rect 1489 13243 1547 13249
rect 1489 13240 1501 13243
rect 1452 13212 1501 13240
rect 1452 13200 1458 13212
rect 1489 13209 1501 13212
rect 1535 13209 1547 13243
rect 1489 13203 1547 13209
rect 6638 13200 6644 13252
rect 6696 13200 6702 13252
rect 15470 13240 15476 13252
rect 8220 13212 15476 13240
rect 1578 13132 1584 13184
rect 1636 13172 1642 13184
rect 8220 13181 8248 13212
rect 15470 13200 15476 13212
rect 15528 13200 15534 13252
rect 2777 13175 2835 13181
rect 2777 13172 2789 13175
rect 1636 13144 2789 13172
rect 1636 13132 1642 13144
rect 2777 13141 2789 13144
rect 2823 13141 2835 13175
rect 2777 13135 2835 13141
rect 8205 13175 8263 13181
rect 8205 13141 8217 13175
rect 8251 13141 8263 13175
rect 8205 13135 8263 13141
rect 920 13082 9844 13104
rect 920 13030 3566 13082
rect 3618 13030 3630 13082
rect 3682 13030 3694 13082
rect 3746 13030 3758 13082
rect 3810 13030 3822 13082
rect 3874 13030 8566 13082
rect 8618 13030 8630 13082
rect 8682 13030 8694 13082
rect 8746 13030 8758 13082
rect 8810 13030 8822 13082
rect 8874 13030 9844 13082
rect 920 13008 9844 13030
rect 8294 12968 8300 12980
rect 8255 12940 8300 12968
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 17310 12968 17316 12980
rect 13872 12940 17316 12968
rect 13872 12928 13878 12940
rect 17310 12928 17316 12940
rect 17368 12928 17374 12980
rect 3510 12860 3516 12912
rect 3568 12860 3574 12912
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 1762 12832 1768 12844
rect 1627 12804 1768 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 2958 12832 2964 12844
rect 2919 12804 2964 12832
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 4430 12832 4436 12844
rect 4391 12804 4436 12832
rect 4430 12792 4436 12804
rect 4488 12792 4494 12844
rect 5258 12792 5264 12844
rect 5316 12832 5322 12844
rect 5353 12835 5411 12841
rect 5353 12832 5365 12835
rect 5316 12804 5365 12832
rect 5316 12792 5322 12804
rect 5353 12801 5365 12804
rect 5399 12801 5411 12835
rect 6546 12832 6552 12844
rect 6507 12804 6552 12832
rect 5353 12795 5411 12801
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 7926 12792 7932 12844
rect 7984 12792 7990 12844
rect 9217 12835 9275 12841
rect 9217 12801 9229 12835
rect 9263 12832 9275 12835
rect 15010 12832 15016 12844
rect 9263 12804 15016 12832
rect 9263 12801 9275 12804
rect 9217 12795 9275 12801
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 5629 12767 5687 12773
rect 5629 12733 5641 12767
rect 5675 12764 5687 12767
rect 5810 12764 5816 12776
rect 5675 12736 5816 12764
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 5810 12724 5816 12736
rect 5868 12724 5874 12776
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 7190 12764 7196 12776
rect 6871 12736 7196 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 13446 12656 13452 12708
rect 13504 12696 13510 12708
rect 15194 12696 15200 12708
rect 13504 12668 15200 12696
rect 13504 12656 13510 12668
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 842 12588 848 12640
rect 900 12628 906 12640
rect 2133 12631 2191 12637
rect 2133 12628 2145 12631
rect 900 12600 2145 12628
rect 900 12588 906 12600
rect 2133 12597 2145 12600
rect 2179 12597 2191 12631
rect 4890 12628 4896 12640
rect 4851 12600 4896 12628
rect 2133 12591 2191 12597
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 9125 12631 9183 12637
rect 9125 12628 9137 12631
rect 7984 12600 9137 12628
rect 7984 12588 7990 12600
rect 9125 12597 9137 12600
rect 9171 12628 9183 12631
rect 9490 12628 9496 12640
rect 9171 12600 9496 12628
rect 9171 12597 9183 12600
rect 9125 12591 9183 12597
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 920 12538 9844 12560
rect 920 12486 2566 12538
rect 2618 12486 2630 12538
rect 2682 12486 2694 12538
rect 2746 12486 2758 12538
rect 2810 12486 2822 12538
rect 2874 12486 7566 12538
rect 7618 12486 7630 12538
rect 7682 12486 7694 12538
rect 7746 12486 7758 12538
rect 7810 12486 7822 12538
rect 7874 12486 9844 12538
rect 13814 12520 13820 12572
rect 13872 12560 13878 12572
rect 15930 12560 15936 12572
rect 13872 12532 15936 12560
rect 13872 12520 13878 12532
rect 15930 12520 15936 12532
rect 15988 12520 15994 12572
rect 920 12464 9844 12486
rect 658 12384 664 12436
rect 716 12424 722 12436
rect 1210 12424 1216 12436
rect 716 12396 1216 12424
rect 716 12384 722 12396
rect 1210 12384 1216 12396
rect 1268 12384 1274 12436
rect 2406 12248 2412 12300
rect 2464 12288 2470 12300
rect 2961 12291 3019 12297
rect 2961 12288 2973 12291
rect 2464 12260 2973 12288
rect 2464 12248 2470 12260
rect 2961 12257 2973 12260
rect 3007 12257 3019 12291
rect 2961 12251 3019 12257
rect 13832 12260 15194 12288
rect 13832 12232 13860 12260
rect 3234 12180 3240 12232
rect 3292 12220 3298 12232
rect 3418 12220 3424 12232
rect 3292 12192 3424 12220
rect 3292 12180 3298 12192
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12220 4031 12223
rect 4062 12220 4068 12232
rect 4019 12192 4068 12220
rect 4019 12189 4031 12192
rect 3973 12183 4031 12189
rect 3050 12152 3056 12164
rect 2530 12124 3056 12152
rect 3050 12112 3056 12124
rect 3108 12112 3114 12164
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 2958 12044 2964 12096
rect 3016 12084 3022 12096
rect 3804 12084 3832 12183
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 4433 12223 4491 12229
rect 4433 12220 4445 12223
rect 4304 12192 4445 12220
rect 4304 12180 4310 12192
rect 4433 12189 4445 12192
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 4706 12180 4712 12232
rect 4764 12220 4770 12232
rect 4801 12223 4859 12229
rect 4801 12220 4813 12223
rect 4764 12192 4813 12220
rect 4764 12180 4770 12192
rect 4801 12189 4813 12192
rect 4847 12189 4859 12223
rect 6270 12220 6276 12232
rect 6231 12192 6276 12220
rect 4801 12183 4859 12189
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7558 12220 7564 12232
rect 7248 12192 7564 12220
rect 7248 12180 7254 12192
rect 7558 12180 7564 12192
rect 7616 12180 7622 12232
rect 8754 12180 8760 12232
rect 8812 12220 8818 12232
rect 8941 12223 8999 12229
rect 8941 12220 8953 12223
rect 8812 12192 8953 12220
rect 8812 12180 8818 12192
rect 8941 12189 8953 12192
rect 8987 12189 8999 12223
rect 8941 12183 8999 12189
rect 12342 12180 12348 12232
rect 12400 12220 12406 12232
rect 12986 12220 12992 12232
rect 12400 12192 12992 12220
rect 12400 12180 12406 12192
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 13814 12180 13820 12232
rect 13872 12180 13878 12232
rect 15010 12180 15016 12232
rect 15068 12220 15074 12232
rect 15166 12220 15194 12260
rect 15838 12220 15844 12232
rect 15068 12192 15844 12220
rect 15068 12180 15074 12192
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 5902 12112 5908 12164
rect 5960 12112 5966 12164
rect 7098 12112 7104 12164
rect 7156 12152 7162 12164
rect 7926 12152 7932 12164
rect 7156 12124 7932 12152
rect 7156 12112 7162 12124
rect 7926 12112 7932 12124
rect 7984 12112 7990 12164
rect 8202 12112 8208 12164
rect 8260 12152 8266 12164
rect 9125 12155 9183 12161
rect 9125 12152 9137 12155
rect 8260 12124 9137 12152
rect 8260 12112 8266 12124
rect 9125 12121 9137 12124
rect 9171 12152 9183 12155
rect 9398 12152 9404 12164
rect 9171 12124 9404 12152
rect 9171 12121 9183 12124
rect 9125 12115 9183 12121
rect 9398 12112 9404 12124
rect 9456 12112 9462 12164
rect 3016 12056 3832 12084
rect 3881 12087 3939 12093
rect 3016 12044 3022 12056
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 4062 12084 4068 12096
rect 3927 12056 4068 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 6546 12044 6552 12096
rect 6604 12084 6610 12096
rect 6733 12087 6791 12093
rect 6733 12084 6745 12087
rect 6604 12056 6745 12084
rect 6604 12044 6610 12056
rect 6733 12053 6745 12056
rect 6779 12053 6791 12087
rect 6733 12047 6791 12053
rect 8113 12087 8171 12093
rect 8113 12053 8125 12087
rect 8159 12084 8171 12087
rect 8294 12084 8300 12096
rect 8159 12056 8300 12084
rect 8159 12053 8171 12056
rect 8113 12047 8171 12053
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 9306 12084 9312 12096
rect 9267 12056 9312 12084
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 920 11994 9844 12016
rect 920 11942 3566 11994
rect 3618 11942 3630 11994
rect 3682 11942 3694 11994
rect 3746 11942 3758 11994
rect 3810 11942 3822 11994
rect 3874 11942 8566 11994
rect 8618 11942 8630 11994
rect 8682 11942 8694 11994
rect 8746 11942 8758 11994
rect 8810 11942 8822 11994
rect 8874 11942 9844 11994
rect 920 11920 9844 11942
rect 13814 11908 13820 11960
rect 13872 11948 13878 11960
rect 15470 11948 15476 11960
rect 13872 11920 15476 11948
rect 13872 11908 13878 11920
rect 15470 11908 15476 11920
rect 15528 11908 15534 11960
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 8113 11883 8171 11889
rect 8113 11880 8125 11883
rect 7616 11852 8125 11880
rect 7616 11840 7622 11852
rect 8113 11849 8125 11852
rect 8159 11849 8171 11883
rect 8113 11843 8171 11849
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 9088 11852 9229 11880
rect 9088 11840 9094 11852
rect 9217 11849 9229 11852
rect 9263 11849 9275 11883
rect 9217 11843 9275 11849
rect 3050 11812 3056 11824
rect 2898 11784 3056 11812
rect 3050 11772 3056 11784
rect 3108 11772 3114 11824
rect 5810 11812 5816 11824
rect 5771 11784 5816 11812
rect 5810 11772 5816 11784
rect 5868 11772 5874 11824
rect 7098 11772 7104 11824
rect 7156 11772 7162 11824
rect 8849 11815 8907 11821
rect 8849 11781 8861 11815
rect 8895 11812 8907 11815
rect 13538 11812 13544 11824
rect 8895 11784 13544 11812
rect 8895 11781 8907 11784
rect 8849 11775 8907 11781
rect 13538 11772 13544 11784
rect 13596 11772 13602 11824
rect 13814 11772 13820 11824
rect 13872 11812 13878 11824
rect 16482 11812 16488 11824
rect 13872 11784 16488 11812
rect 13872 11772 13878 11784
rect 16482 11772 16488 11784
rect 16540 11772 16546 11824
rect 8754 11744 8760 11756
rect 8715 11716 8760 11744
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 8938 11704 8944 11756
rect 8996 11744 9002 11756
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8996 11716 9045 11744
rect 8996 11704 9002 11716
rect 9033 11713 9045 11716
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 3234 11636 3240 11688
rect 3292 11676 3298 11688
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 3292 11648 3341 11676
rect 3292 11636 3298 11648
rect 3329 11645 3341 11648
rect 3375 11645 3387 11679
rect 3602 11676 3608 11688
rect 3563 11648 3608 11676
rect 3329 11639 3387 11645
rect 3602 11636 3608 11648
rect 3660 11636 3666 11688
rect 4154 11676 4160 11688
rect 4115 11648 4160 11676
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 6362 11676 6368 11688
rect 6323 11648 6368 11676
rect 6362 11636 6368 11648
rect 6420 11636 6426 11688
rect 6638 11676 6644 11688
rect 6599 11648 6644 11676
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 1854 11540 1860 11552
rect 1815 11512 1860 11540
rect 1854 11500 1860 11512
rect 1912 11500 1918 11552
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 7566 11450
rect 7618 11398 7630 11450
rect 7682 11398 7694 11450
rect 7746 11398 7758 11450
rect 7810 11398 7822 11450
rect 7874 11398 9844 11450
rect 13538 11432 13544 11484
rect 13596 11472 13602 11484
rect 15654 11472 15660 11484
rect 13596 11444 15660 11472
rect 13596 11432 13602 11444
rect 15654 11432 15660 11444
rect 15712 11432 15718 11484
rect 920 11376 9844 11398
rect 2130 11336 2136 11348
rect 2091 11308 2136 11336
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2682 11200 2688 11212
rect 2643 11172 2688 11200
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4614 11200 4620 11212
rect 4479 11172 4620 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 1854 11132 1860 11144
rect 1627 11104 1860 11132
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 1854 11092 1860 11104
rect 1912 11132 1918 11144
rect 1912 11104 2774 11132
rect 1912 11092 1918 11104
rect 2746 10996 2774 11104
rect 5810 11092 5816 11144
rect 5868 11132 5874 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 5868 11104 8033 11132
rect 5868 11092 5874 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8536 11104 8953 11132
rect 8536 11092 8542 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 3234 11064 3240 11076
rect 3195 11036 3240 11064
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 5534 11064 5540 11076
rect 5495 11036 5540 11064
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 7190 11064 7196 11076
rect 7151 11036 7196 11064
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 7466 11024 7472 11076
rect 7524 11064 7530 11076
rect 7653 11067 7711 11073
rect 7653 11064 7665 11067
rect 7524 11036 7665 11064
rect 7524 11024 7530 11036
rect 7653 11033 7665 11036
rect 7699 11033 7711 11067
rect 7837 11067 7895 11073
rect 7837 11064 7849 11067
rect 7653 11027 7711 11033
rect 7760 11036 7849 11064
rect 4062 10996 4068 11008
rect 2746 10968 4068 10996
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 4985 10999 5043 11005
rect 4985 10965 4997 10999
rect 5031 10996 5043 10999
rect 5166 10996 5172 11008
rect 5031 10968 5172 10996
rect 5031 10965 5043 10968
rect 4985 10959 5043 10965
rect 5166 10956 5172 10968
rect 5224 10956 5230 11008
rect 5626 10956 5632 11008
rect 5684 10996 5690 11008
rect 7760 10996 7788 11036
rect 7837 11033 7849 11036
rect 7883 11064 7895 11067
rect 8202 11064 8208 11076
rect 7883 11036 8208 11064
rect 7883 11033 7895 11036
rect 7837 11027 7895 11033
rect 8202 11024 8208 11036
rect 8260 11024 8266 11076
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 18138 11064 18144 11076
rect 14884 11036 18144 11064
rect 14884 11024 14890 11036
rect 18138 11024 18144 11036
rect 18196 11024 18202 11076
rect 5684 10968 7788 10996
rect 9125 10999 9183 11005
rect 5684 10956 5690 10968
rect 9125 10965 9137 10999
rect 9171 10996 9183 10999
rect 14090 10996 14096 11008
rect 9171 10968 14096 10996
rect 9171 10965 9183 10968
rect 9125 10959 9183 10965
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 920 10906 9844 10928
rect 920 10854 3566 10906
rect 3618 10854 3630 10906
rect 3682 10854 3694 10906
rect 3746 10854 3758 10906
rect 3810 10854 3822 10906
rect 3874 10854 8566 10906
rect 8618 10854 8630 10906
rect 8682 10854 8694 10906
rect 8746 10854 8758 10906
rect 8810 10854 8822 10906
rect 8874 10854 9844 10906
rect 920 10832 9844 10854
rect 4798 10792 4804 10804
rect 4759 10764 4804 10792
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 3878 10684 3884 10736
rect 3936 10684 3942 10736
rect 5445 10727 5503 10733
rect 5445 10693 5457 10727
rect 5491 10724 5503 10727
rect 5718 10724 5724 10736
rect 5491 10696 5724 10724
rect 5491 10693 5503 10696
rect 5445 10687 5503 10693
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 7190 10684 7196 10736
rect 7248 10684 7254 10736
rect 1489 10659 1547 10665
rect 1489 10625 1501 10659
rect 1535 10656 1547 10659
rect 1670 10656 1676 10668
rect 1535 10628 1676 10656
rect 1535 10625 1547 10628
rect 1489 10619 1547 10625
rect 1670 10616 1676 10628
rect 1728 10616 1734 10668
rect 2130 10616 2136 10668
rect 2188 10656 2194 10668
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2188 10628 2881 10656
rect 2188 10616 2194 10628
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 4338 10656 4344 10668
rect 4299 10628 4344 10656
rect 2869 10619 2927 10625
rect 4338 10616 4344 10628
rect 4396 10616 4402 10668
rect 5626 10656 5632 10668
rect 5587 10628 5632 10656
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 6178 10616 6184 10668
rect 6236 10656 6242 10668
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6236 10628 6837 10656
rect 6236 10616 6242 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 8294 10656 8300 10668
rect 8255 10628 8300 10656
rect 6825 10619 6883 10625
rect 8294 10616 8300 10628
rect 8352 10616 8358 10668
rect 8386 10616 8392 10668
rect 8444 10656 8450 10668
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 8444 10628 9137 10656
rect 8444 10616 8450 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 2498 10588 2504 10600
rect 2459 10560 2504 10588
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10588 8723 10591
rect 9217 10591 9275 10597
rect 9217 10588 9229 10591
rect 8711 10560 9229 10588
rect 8711 10557 8723 10560
rect 8665 10551 8723 10557
rect 9217 10557 9229 10560
rect 9263 10557 9275 10591
rect 9217 10551 9275 10557
rect 5813 10523 5871 10529
rect 5813 10489 5825 10523
rect 5859 10520 5871 10523
rect 6730 10520 6736 10532
rect 5859 10492 6736 10520
rect 5859 10489 5871 10492
rect 5813 10483 5871 10489
rect 6730 10480 6736 10492
rect 6788 10480 6794 10532
rect 13814 10480 13820 10532
rect 13872 10520 13878 10532
rect 16942 10520 16948 10532
rect 13872 10492 16948 10520
rect 13872 10480 13878 10492
rect 16942 10480 16948 10492
rect 17000 10480 17006 10532
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 6328 10424 6377 10452
rect 6328 10412 6334 10424
rect 6365 10421 6377 10424
rect 6411 10421 6423 10455
rect 6365 10415 6423 10421
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 7566 10362
rect 7618 10310 7630 10362
rect 7682 10310 7694 10362
rect 7746 10310 7758 10362
rect 7810 10310 7822 10362
rect 7874 10310 9844 10362
rect 920 10288 9844 10310
rect 13814 10276 13820 10328
rect 13872 10316 13878 10328
rect 18414 10316 18420 10328
rect 13872 10288 18420 10316
rect 13872 10276 13878 10288
rect 18414 10276 18420 10288
rect 18472 10276 18478 10328
rect 2130 10248 2136 10260
rect 2091 10220 2136 10248
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 8938 10248 8944 10260
rect 8899 10220 8944 10248
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9122 10248 9128 10260
rect 9083 10220 9128 10248
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 13722 10140 13728 10192
rect 13780 10180 13786 10192
rect 18414 10180 18420 10192
rect 13780 10152 18420 10180
rect 13780 10140 13786 10152
rect 18414 10140 18420 10152
rect 18472 10140 18478 10192
rect 1486 10112 1492 10124
rect 1447 10084 1492 10112
rect 1486 10072 1492 10084
rect 1544 10072 1550 10124
rect 2314 10072 2320 10124
rect 2372 10112 2378 10124
rect 2593 10115 2651 10121
rect 2593 10112 2605 10115
rect 2372 10084 2605 10112
rect 2372 10072 2378 10084
rect 2593 10081 2605 10084
rect 2639 10081 2651 10115
rect 4062 10112 4068 10124
rect 4023 10084 4068 10112
rect 2593 10075 2651 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10112 8355 10115
rect 9674 10112 9680 10124
rect 8343 10084 9680 10112
rect 8343 10081 8355 10084
rect 8297 10075 8355 10081
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 15562 10112 15568 10124
rect 10560 10084 15568 10112
rect 10560 10072 10566 10084
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 3418 10004 3424 10056
rect 3476 10044 3482 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3476 10016 3801 10044
rect 3476 10004 3482 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 5994 10044 6000 10056
rect 5955 10016 6000 10044
rect 3789 10007 3847 10013
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6362 10044 6368 10056
rect 6323 10016 6368 10044
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 8110 10044 8116 10056
rect 7883 10016 8116 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 5442 9976 5448 9988
rect 5290 9948 5448 9976
rect 5442 9936 5448 9948
rect 5500 9936 5506 9988
rect 7006 9936 7012 9988
rect 7064 9936 7070 9988
rect 9306 9976 9312 9988
rect 9267 9948 9312 9976
rect 9306 9936 9312 9948
rect 9364 9936 9370 9988
rect 3234 9908 3240 9920
rect 3195 9880 3240 9908
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 3878 9868 3884 9920
rect 3936 9908 3942 9920
rect 4062 9908 4068 9920
rect 3936 9880 4068 9908
rect 3936 9868 3942 9880
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 5537 9911 5595 9917
rect 5537 9877 5549 9911
rect 5583 9908 5595 9911
rect 6638 9908 6644 9920
rect 5583 9880 6644 9908
rect 5583 9877 5595 9880
rect 5537 9871 5595 9877
rect 6638 9868 6644 9880
rect 6696 9908 6702 9920
rect 6822 9908 6828 9920
rect 6696 9880 6828 9908
rect 6696 9868 6702 9880
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 8018 9908 8024 9920
rect 7979 9880 8024 9908
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 9109 9911 9167 9917
rect 9109 9908 9121 9911
rect 8352 9880 9121 9908
rect 8352 9868 8358 9880
rect 9109 9877 9121 9880
rect 9155 9908 9167 9911
rect 13906 9908 13912 9920
rect 9155 9880 13912 9908
rect 9155 9877 9167 9880
rect 9109 9871 9167 9877
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 14090 9868 14096 9920
rect 14148 9908 14154 9920
rect 15470 9908 15476 9920
rect 14148 9880 15476 9908
rect 14148 9868 14154 9880
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 920 9818 9844 9840
rect 920 9766 3566 9818
rect 3618 9766 3630 9818
rect 3682 9766 3694 9818
rect 3746 9766 3758 9818
rect 3810 9766 3822 9818
rect 3874 9766 8566 9818
rect 8618 9766 8630 9818
rect 8682 9766 8694 9818
rect 8746 9766 8758 9818
rect 8810 9766 8822 9818
rect 8874 9766 9844 9818
rect 920 9744 9844 9766
rect 9306 9704 9312 9716
rect 7208 9676 9312 9704
rect 4614 9596 4620 9648
rect 4672 9596 4678 9648
rect 7208 9636 7236 9676
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 7374 9636 7380 9648
rect 6472 9608 7236 9636
rect 7335 9608 7380 9636
rect 6472 9580 6500 9608
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 9125 9639 9183 9645
rect 9125 9605 9137 9639
rect 9171 9636 9183 9639
rect 15286 9636 15292 9648
rect 9171 9608 15292 9636
rect 9171 9605 9183 9608
rect 9125 9599 9183 9605
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 3053 9571 3111 9577
rect 3053 9537 3065 9571
rect 3099 9568 3111 9571
rect 3234 9568 3240 9580
rect 3099 9540 3240 9568
rect 3099 9537 3111 9540
rect 3053 9531 3111 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9568 3571 9571
rect 3970 9568 3976 9580
rect 3559 9540 3976 9568
rect 3559 9537 3571 9540
rect 3513 9531 3571 9537
rect 3970 9528 3976 9540
rect 4028 9528 4034 9580
rect 5350 9568 5356 9580
rect 5311 9540 5356 9568
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 6454 9568 6460 9580
rect 6415 9540 6460 9568
rect 6454 9528 6460 9540
rect 6512 9528 6518 9580
rect 1489 9503 1547 9509
rect 1489 9469 1501 9503
rect 1535 9500 1547 9503
rect 2130 9500 2136 9512
rect 1535 9472 2136 9500
rect 1535 9469 1547 9472
rect 1489 9463 1547 9469
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 2682 9500 2688 9512
rect 2643 9472 2688 9500
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3016 9472 3893 9500
rect 3016 9460 3022 9472
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 5810 9500 5816 9512
rect 5771 9472 5816 9500
rect 3881 9463 3939 9469
rect 5810 9460 5816 9472
rect 5868 9460 5874 9512
rect 13170 9460 13176 9512
rect 13228 9500 13234 9512
rect 18046 9500 18052 9512
rect 13228 9472 18052 9500
rect 13228 9460 13234 9472
rect 18046 9460 18052 9472
rect 18104 9460 18110 9512
rect 4982 9392 4988 9444
rect 5040 9432 5046 9444
rect 5040 9404 6592 9432
rect 5040 9392 5046 9404
rect 6564 9373 6592 9404
rect 6549 9367 6607 9373
rect 6549 9333 6561 9367
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 6917 9367 6975 9373
rect 6917 9333 6929 9367
rect 6963 9364 6975 9367
rect 9030 9364 9036 9376
rect 6963 9336 9036 9364
rect 6963 9333 6975 9336
rect 6917 9327 6975 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 7566 9274
rect 7618 9222 7630 9274
rect 7682 9222 7694 9274
rect 7746 9222 7758 9274
rect 7810 9222 7822 9274
rect 7874 9222 9844 9274
rect 920 9200 9844 9222
rect 13814 9188 13820 9240
rect 13872 9228 13878 9240
rect 15470 9228 15476 9240
rect 13872 9200 15476 9228
rect 13872 9188 13878 9200
rect 15470 9188 15476 9200
rect 15528 9188 15534 9240
rect 4706 9160 4712 9172
rect 4667 9132 4712 9160
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 1486 9052 1492 9104
rect 1544 9052 1550 9104
rect 13814 9052 13820 9104
rect 13872 9092 13878 9104
rect 15746 9092 15752 9104
rect 13872 9064 15752 9092
rect 13872 9052 13878 9064
rect 15746 9052 15752 9064
rect 15804 9052 15810 9104
rect 1504 9024 1532 9052
rect 1765 9027 1823 9033
rect 1765 9024 1777 9027
rect 1504 8996 1777 9024
rect 1765 8993 1777 8996
rect 1811 8993 1823 9027
rect 1765 8987 1823 8993
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 3200 8996 4077 9024
rect 3200 8984 3206 8996
rect 4065 8993 4077 8996
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7653 9027 7711 9033
rect 7653 9024 7665 9027
rect 7156 8996 7665 9024
rect 7156 8984 7162 8996
rect 7653 8993 7665 8996
rect 7699 8993 7711 9027
rect 7653 8987 7711 8993
rect 14274 8984 14280 9036
rect 14332 9024 14338 9036
rect 15378 9024 15384 9036
rect 14332 8996 15384 9024
rect 14332 8984 14338 8996
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 1486 8956 1492 8968
rect 1447 8928 1492 8956
rect 1486 8916 1492 8928
rect 1544 8916 1550 8968
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 5261 8959 5319 8965
rect 5261 8956 5273 8959
rect 4212 8928 5273 8956
rect 4212 8916 4218 8928
rect 5261 8925 5273 8928
rect 5307 8956 5319 8959
rect 5442 8956 5448 8968
rect 5307 8928 5448 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 7282 8916 7288 8968
rect 7340 8956 7346 8968
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 7340 8928 7481 8956
rect 7340 8916 7346 8928
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 9030 8956 9036 8968
rect 8991 8928 9036 8956
rect 7469 8919 7527 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 13078 8916 13084 8968
rect 13136 8956 13142 8968
rect 17678 8956 17684 8968
rect 13136 8928 17684 8956
rect 13136 8916 13142 8928
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 2314 8848 2320 8900
rect 2372 8848 2378 8900
rect 15378 8848 15384 8900
rect 15436 8888 15442 8900
rect 15930 8888 15936 8900
rect 15436 8860 15936 8888
rect 15436 8848 15442 8860
rect 15930 8848 15936 8860
rect 15988 8848 15994 8900
rect 1762 8780 1768 8832
rect 1820 8820 1826 8832
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 1820 8792 3249 8820
rect 1820 8780 1826 8792
rect 3237 8789 3249 8792
rect 3283 8789 3295 8823
rect 3237 8783 3295 8789
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 4948 8792 6561 8820
rect 4948 8780 4954 8792
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 9122 8820 9128 8832
rect 9083 8792 9128 8820
rect 6549 8783 6607 8789
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 920 8730 9844 8752
rect 920 8678 3566 8730
rect 3618 8678 3630 8730
rect 3682 8678 3694 8730
rect 3746 8678 3758 8730
rect 3810 8678 3822 8730
rect 3874 8678 8566 8730
rect 8618 8678 8630 8730
rect 8682 8678 8694 8730
rect 8746 8678 8758 8730
rect 8810 8678 8822 8730
rect 8874 8678 9844 8730
rect 920 8656 9844 8678
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 5040 8588 5089 8616
rect 5040 8576 5046 8588
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 5626 8616 5632 8628
rect 5587 8588 5632 8616
rect 5077 8579 5135 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 6362 8616 6368 8628
rect 6323 8588 6368 8616
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 3510 8508 3516 8560
rect 3568 8508 3574 8560
rect 9122 8548 9128 8560
rect 9083 8520 9128 8548
rect 9122 8508 9128 8520
rect 9180 8508 9186 8560
rect 1762 8480 1768 8492
rect 1723 8452 1768 8480
rect 1762 8440 1768 8452
rect 1820 8440 1826 8492
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 3145 8483 3203 8489
rect 3145 8480 3157 8483
rect 2363 8452 3157 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 3145 8449 3157 8452
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 4430 8440 4436 8492
rect 4488 8480 4494 8492
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 4488 8452 4629 8480
rect 4488 8440 4494 8452
rect 4617 8449 4629 8452
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 5994 8480 6000 8492
rect 5859 8452 6000 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6914 8480 6920 8492
rect 6875 8452 6920 8480
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 15194 8480 15200 8492
rect 11296 8452 15200 8480
rect 11296 8440 11302 8452
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 8202 8412 8208 8424
rect 2832 8384 2877 8412
rect 8163 8384 8208 8412
rect 2832 8372 2838 8384
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8412 9367 8415
rect 9582 8412 9588 8424
rect 9355 8384 9588 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 6454 8304 6460 8356
rect 6512 8344 6518 8356
rect 7098 8344 7104 8356
rect 6512 8316 7104 8344
rect 6512 8304 6518 8316
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 13538 8304 13544 8356
rect 13596 8344 13602 8356
rect 18506 8344 18512 8356
rect 13596 8316 18512 8344
rect 13596 8304 13602 8316
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 16022 8276 16028 8288
rect 13320 8248 16028 8276
rect 13320 8236 13326 8248
rect 16022 8236 16028 8248
rect 16080 8236 16086 8288
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 7566 8186
rect 7618 8134 7630 8186
rect 7682 8134 7694 8186
rect 7746 8134 7758 8186
rect 7810 8134 7822 8186
rect 7874 8134 9844 8186
rect 920 8112 9844 8134
rect 3878 7936 3884 7948
rect 3839 7908 3884 7936
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 1394 7828 1400 7880
rect 1452 7868 1458 7880
rect 1489 7871 1547 7877
rect 1489 7868 1501 7871
rect 1452 7840 1501 7868
rect 1452 7828 1458 7840
rect 1489 7837 1501 7840
rect 1535 7837 1547 7871
rect 1489 7831 1547 7837
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7374 7868 7380 7880
rect 7055 7840 7380 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 8018 7868 8024 7880
rect 7979 7840 8024 7868
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8536 7840 8953 7868
rect 8536 7828 8542 7840
rect 8941 7837 8953 7840
rect 8987 7868 8999 7871
rect 9490 7868 9496 7880
rect 8987 7840 9496 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 3234 7800 3240 7812
rect 3195 7772 3240 7800
rect 3234 7760 3240 7772
rect 3292 7760 3298 7812
rect 5258 7800 5264 7812
rect 5219 7772 5264 7800
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 9125 7803 9183 7809
rect 9125 7769 9137 7803
rect 9171 7800 9183 7803
rect 9214 7800 9220 7812
rect 9171 7772 9220 7800
rect 9171 7769 9183 7772
rect 9125 7763 9183 7769
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 4430 7732 4436 7744
rect 4391 7704 4436 7732
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7469 7735 7527 7741
rect 7469 7732 7481 7735
rect 7064 7704 7481 7732
rect 7064 7692 7070 7704
rect 7469 7701 7481 7704
rect 7515 7701 7527 7735
rect 7469 7695 7527 7701
rect 9309 7735 9367 7741
rect 9309 7701 9321 7735
rect 9355 7732 9367 7735
rect 9858 7732 9864 7744
rect 9355 7704 9864 7732
rect 9355 7701 9367 7704
rect 9309 7695 9367 7701
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 920 7642 9844 7664
rect 920 7590 3566 7642
rect 3618 7590 3630 7642
rect 3682 7590 3694 7642
rect 3746 7590 3758 7642
rect 3810 7590 3822 7642
rect 3874 7590 8566 7642
rect 8618 7590 8630 7642
rect 8682 7590 8694 7642
rect 8746 7590 8758 7642
rect 8810 7590 8822 7642
rect 8874 7590 9844 7642
rect 11330 7624 11336 7676
rect 11388 7664 11394 7676
rect 15838 7664 15844 7676
rect 11388 7636 15844 7664
rect 11388 7624 11394 7636
rect 15838 7624 15844 7636
rect 15896 7624 15902 7676
rect 920 7568 9844 7590
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 5684 7500 5825 7528
rect 5684 7488 5690 7500
rect 5813 7497 5825 7500
rect 5859 7528 5871 7531
rect 8018 7528 8024 7540
rect 5859 7500 8024 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 9122 7528 9128 7540
rect 9083 7500 9128 7528
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 1857 7463 1915 7469
rect 1857 7460 1869 7463
rect 1544 7432 1869 7460
rect 1544 7420 1550 7432
rect 1857 7429 1869 7432
rect 1903 7460 1915 7463
rect 3418 7460 3424 7472
rect 1903 7432 3424 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 3418 7420 3424 7432
rect 3476 7420 3482 7472
rect 3605 7463 3663 7469
rect 3605 7429 3617 7463
rect 3651 7460 3663 7463
rect 4062 7460 4068 7472
rect 3651 7432 4068 7460
rect 3651 7429 3663 7432
rect 3605 7423 3663 7429
rect 4062 7420 4068 7432
rect 4120 7420 4126 7472
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 4341 7463 4399 7469
rect 4341 7460 4353 7463
rect 4304 7432 4353 7460
rect 4304 7420 4310 7432
rect 4341 7429 4353 7432
rect 4387 7429 4399 7463
rect 4341 7423 4399 7429
rect 4798 7420 4804 7472
rect 4856 7420 4862 7472
rect 7098 7420 7104 7472
rect 7156 7420 7162 7472
rect 13814 7420 13820 7472
rect 13872 7460 13878 7472
rect 18046 7460 18052 7472
rect 13872 7432 18052 7460
rect 13872 7420 13878 7432
rect 18046 7420 18052 7432
rect 18104 7420 18110 7472
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 8076 7364 8217 7392
rect 8076 7352 8082 7364
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 9306 7392 9312 7404
rect 9267 7364 9312 7392
rect 8205 7355 8263 7361
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 3418 7284 3424 7336
rect 3476 7324 3482 7336
rect 4065 7327 4123 7333
rect 4065 7324 4077 7327
rect 3476 7296 4077 7324
rect 3476 7284 3482 7296
rect 4065 7293 4077 7296
rect 4111 7293 4123 7327
rect 6362 7324 6368 7336
rect 6323 7296 6368 7324
rect 4065 7287 4123 7293
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 6733 7327 6791 7333
rect 6733 7293 6745 7327
rect 6779 7324 6791 7327
rect 6914 7324 6920 7336
rect 6779 7296 6920 7324
rect 6779 7293 6791 7296
rect 6733 7287 6791 7293
rect 6914 7284 6920 7296
rect 6972 7284 6978 7336
rect 8665 7191 8723 7197
rect 8665 7157 8677 7191
rect 8711 7188 8723 7191
rect 8938 7188 8944 7200
rect 8711 7160 8944 7188
rect 8711 7157 8723 7160
rect 8665 7151 8723 7157
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 7566 7098
rect 7618 7046 7630 7098
rect 7682 7046 7694 7098
rect 7746 7046 7758 7098
rect 7810 7046 7822 7098
rect 7874 7046 9844 7098
rect 920 7024 9844 7046
rect 4246 6916 4252 6928
rect 4080 6888 4252 6916
rect 1486 6848 1492 6860
rect 1447 6820 1492 6848
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 1762 6848 1768 6860
rect 1723 6820 1768 6848
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 2314 6808 2320 6860
rect 2372 6848 2378 6860
rect 3881 6851 3939 6857
rect 2372 6820 2912 6848
rect 2372 6808 2378 6820
rect 198 6740 204 6792
rect 256 6780 262 6792
rect 1394 6780 1400 6792
rect 256 6752 1400 6780
rect 256 6740 262 6752
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 2884 6780 2912 6820
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 4080 6848 4108 6888
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 4798 6848 4804 6860
rect 3927 6820 4108 6848
rect 4356 6820 4804 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 4356 6780 4384 6820
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 2884 6766 4384 6780
rect 2898 6752 4384 6766
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 6086 6780 6092 6792
rect 5684 6752 5729 6780
rect 6047 6752 6092 6780
rect 5684 6740 5690 6752
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 6454 6780 6460 6792
rect 6415 6752 6460 6780
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7524 6752 7941 6780
rect 7524 6740 7530 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6780 8999 6783
rect 9030 6780 9036 6792
rect 8987 6752 9036 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 9030 6740 9036 6752
rect 9088 6740 9094 6792
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9214 6780 9220 6792
rect 9171 6752 9220 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 15654 6780 15660 6792
rect 13872 6752 15660 6780
rect 13872 6740 13878 6752
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 4798 6672 4804 6724
rect 4856 6672 4862 6724
rect 5353 6715 5411 6721
rect 5353 6681 5365 6715
rect 5399 6712 5411 6715
rect 5399 6684 5580 6712
rect 5399 6681 5411 6684
rect 5353 6675 5411 6681
rect 5552 6656 5580 6684
rect 7098 6672 7104 6724
rect 7156 6672 7162 6724
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 3237 6647 3295 6653
rect 3237 6644 3249 6647
rect 3200 6616 3249 6644
rect 3200 6604 3206 6616
rect 3237 6613 3249 6616
rect 3283 6613 3295 6647
rect 3237 6607 3295 6613
rect 5534 6604 5540 6656
rect 5592 6604 5598 6656
rect 8389 6647 8447 6653
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 8478 6644 8484 6656
rect 8435 6616 8484 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 9306 6644 9312 6656
rect 9267 6616 9312 6644
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 920 6554 9844 6576
rect 920 6502 3566 6554
rect 3618 6502 3630 6554
rect 3682 6502 3694 6554
rect 3746 6502 3758 6554
rect 3810 6502 3822 6554
rect 3874 6502 8566 6554
rect 8618 6502 8630 6554
rect 8682 6502 8694 6554
rect 8746 6502 8758 6554
rect 8810 6502 8822 6554
rect 8874 6502 9844 6554
rect 920 6480 9844 6502
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 2682 6440 2688 6452
rect 2363 6412 2688 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 2682 6400 2688 6412
rect 2740 6400 2746 6452
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 3237 6443 3295 6449
rect 3237 6440 3249 6443
rect 3108 6412 3249 6440
rect 3108 6400 3114 6412
rect 3237 6409 3249 6412
rect 3283 6409 3295 6443
rect 3237 6403 3295 6409
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 5626 6440 5632 6452
rect 3476 6412 5632 6440
rect 3476 6400 3482 6412
rect 4798 6372 4804 6384
rect 4278 6344 4804 6372
rect 4798 6332 4804 6344
rect 4856 6332 4862 6384
rect 5000 6313 5028 6412
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 7374 6332 7380 6384
rect 7432 6332 7438 6384
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 6270 6304 6276 6316
rect 5859 6276 6276 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 7006 6304 7012 6316
rect 6963 6276 7012 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6304 8447 6307
rect 9490 6304 9496 6316
rect 8435 6276 9496 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 1765 6239 1823 6245
rect 1765 6205 1777 6239
rect 1811 6236 1823 6239
rect 3142 6236 3148 6248
rect 1811 6208 3148 6236
rect 1811 6205 1823 6208
rect 1765 6199 1823 6205
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 5442 6236 5448 6248
rect 4755 6208 5448 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 6549 6239 6607 6245
rect 6549 6205 6561 6239
rect 6595 6236 6607 6239
rect 6822 6236 6828 6248
rect 6595 6208 6828 6236
rect 6595 6205 6607 6208
rect 6549 6199 6607 6205
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 17908 6128 17914 6180
rect 17966 6168 17972 6180
rect 18598 6168 18604 6180
rect 17966 6140 18604 6168
rect 17966 6128 17972 6140
rect 18598 6128 18604 6140
rect 18656 6128 18662 6180
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 8110 6100 8116 6112
rect 5675 6072 8116 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8849 6103 8907 6109
rect 8849 6069 8861 6103
rect 8895 6100 8907 6103
rect 9122 6100 9128 6112
rect 8895 6072 9128 6100
rect 8895 6069 8907 6072
rect 8849 6063 8907 6069
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 7566 6010
rect 7618 5958 7630 6010
rect 7682 5958 7694 6010
rect 7746 5958 7758 6010
rect 7810 5958 7822 6010
rect 7874 5958 9844 6010
rect 920 5936 9844 5958
rect 1765 5899 1823 5905
rect 1765 5865 1777 5899
rect 1811 5896 1823 5899
rect 2222 5896 2228 5908
rect 1811 5868 2228 5896
rect 1811 5865 1823 5868
rect 1765 5859 1823 5865
rect 2222 5856 2228 5868
rect 2280 5856 2286 5908
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 3053 5899 3111 5905
rect 3053 5896 3065 5899
rect 3016 5868 3065 5896
rect 3016 5856 3022 5868
rect 3053 5865 3065 5868
rect 3099 5865 3111 5899
rect 5534 5896 5540 5908
rect 5495 5868 5540 5896
rect 3053 5859 3111 5865
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 6972 5868 7021 5896
rect 6972 5856 6978 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 8294 5896 8300 5908
rect 8255 5868 8300 5896
rect 7009 5859 7067 5865
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 382 5788 388 5840
rect 440 5828 446 5840
rect 2682 5828 2688 5840
rect 440 5800 2688 5828
rect 440 5788 446 5800
rect 2682 5788 2688 5800
rect 2740 5788 2746 5840
rect 3418 5720 3424 5772
rect 3476 5760 3482 5772
rect 3789 5763 3847 5769
rect 3789 5760 3801 5763
rect 3476 5732 3801 5760
rect 3476 5720 3482 5732
rect 3789 5729 3801 5732
rect 3835 5729 3847 5763
rect 3789 5723 3847 5729
rect 4798 5720 4804 5772
rect 4856 5760 4862 5772
rect 5552 5760 5580 5856
rect 6546 5788 6552 5840
rect 6604 5828 6610 5840
rect 7561 5831 7619 5837
rect 7561 5828 7573 5831
rect 6604 5800 7573 5828
rect 6604 5788 6610 5800
rect 7561 5797 7573 5800
rect 7607 5828 7619 5831
rect 9214 5828 9220 5840
rect 7607 5800 9220 5828
rect 7607 5797 7619 5800
rect 7561 5791 7619 5797
rect 9214 5788 9220 5800
rect 9272 5788 9278 5840
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 15562 5828 15568 5840
rect 13872 5800 15568 5828
rect 13872 5788 13878 5800
rect 15562 5788 15568 5800
rect 15620 5788 15626 5840
rect 6365 5763 6423 5769
rect 6365 5760 6377 5763
rect 4856 5732 5212 5760
rect 5552 5732 6377 5760
rect 4856 5720 4862 5732
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 2498 5692 2504 5704
rect 2459 5664 2504 5692
rect 2498 5652 2504 5664
rect 2556 5652 2562 5704
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3510 5692 3516 5704
rect 3283 5664 3516 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 5184 5692 5212 5732
rect 6365 5729 6377 5732
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 6564 5692 6592 5788
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 9030 5760 9036 5772
rect 8168 5732 9036 5760
rect 8168 5720 8174 5732
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 19058 5720 19064 5772
rect 19116 5720 19122 5772
rect 7742 5692 7748 5704
rect 5184 5678 6592 5692
rect 5198 5664 6592 5678
rect 7703 5664 7748 5692
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 9214 5692 9220 5704
rect 9175 5664 9220 5692
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 19076 5636 19104 5720
rect 1397 5627 1455 5633
rect 1397 5593 1409 5627
rect 1443 5624 1455 5627
rect 1670 5624 1676 5636
rect 1443 5596 1676 5624
rect 1443 5593 1455 5596
rect 1397 5587 1455 5593
rect 1670 5584 1676 5596
rect 1728 5584 1734 5636
rect 3142 5584 3148 5636
rect 3200 5624 3206 5636
rect 4065 5627 4123 5633
rect 4065 5624 4077 5627
rect 3200 5596 4077 5624
rect 3200 5584 3206 5596
rect 4065 5593 4077 5596
rect 4111 5593 4123 5627
rect 4065 5587 4123 5593
rect 7926 5584 7932 5636
rect 7984 5624 7990 5636
rect 8846 5624 8852 5636
rect 7984 5596 8852 5624
rect 7984 5584 7990 5596
rect 8846 5584 8852 5596
rect 8904 5624 8910 5636
rect 8941 5627 8999 5633
rect 8941 5624 8953 5627
rect 8904 5596 8953 5624
rect 8904 5584 8910 5596
rect 8941 5593 8953 5596
rect 8987 5593 8999 5627
rect 8941 5587 8999 5593
rect 9125 5627 9183 5633
rect 9125 5593 9137 5627
rect 9171 5624 9183 5627
rect 10042 5624 10048 5636
rect 9171 5596 10048 5624
rect 9171 5593 9183 5596
rect 9125 5587 9183 5593
rect 10042 5584 10048 5596
rect 10100 5624 10106 5636
rect 13814 5624 13820 5636
rect 10100 5596 13820 5624
rect 10100 5584 10106 5596
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 19058 5584 19064 5636
rect 19116 5584 19122 5636
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5556 2375 5559
rect 2682 5556 2688 5568
rect 2363 5528 2688 5556
rect 2363 5525 2375 5528
rect 2317 5519 2375 5525
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 9030 5556 9036 5568
rect 8991 5528 9036 5556
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 13722 5516 13728 5568
rect 13780 5556 13786 5568
rect 14182 5556 14188 5568
rect 13780 5528 14188 5556
rect 13780 5516 13786 5528
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 920 5466 9844 5488
rect 920 5414 3566 5466
rect 3618 5414 3630 5466
rect 3682 5414 3694 5466
rect 3746 5414 3758 5466
rect 3810 5414 3822 5466
rect 3874 5414 8566 5466
rect 8618 5414 8630 5466
rect 8682 5414 8694 5466
rect 8746 5414 8758 5466
rect 8810 5414 8822 5466
rect 8874 5414 9844 5466
rect 920 5392 9844 5414
rect 106 5312 112 5364
rect 164 5352 170 5364
rect 2498 5352 2504 5364
rect 164 5324 2504 5352
rect 164 5312 170 5324
rect 2498 5312 2504 5324
rect 2556 5312 2562 5364
rect 4062 5352 4068 5364
rect 4023 5324 4068 5352
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 5813 5355 5871 5361
rect 5813 5321 5825 5355
rect 5859 5352 5871 5355
rect 6454 5352 6460 5364
rect 5859 5324 6460 5352
rect 5859 5321 5871 5324
rect 5813 5315 5871 5321
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 7285 5355 7343 5361
rect 7285 5352 7297 5355
rect 6972 5324 7297 5352
rect 6972 5312 6978 5324
rect 7285 5321 7297 5324
rect 7331 5321 7343 5355
rect 7285 5315 7343 5321
rect 8202 5312 8208 5364
rect 8260 5352 8266 5364
rect 9950 5352 9956 5364
rect 8260 5324 9956 5352
rect 8260 5312 8266 5324
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 658 5244 664 5296
rect 716 5284 722 5296
rect 2314 5284 2320 5296
rect 716 5256 2320 5284
rect 716 5244 722 5256
rect 2314 5244 2320 5256
rect 2372 5244 2378 5296
rect 4890 5244 4896 5296
rect 4948 5284 4954 5296
rect 6365 5287 6423 5293
rect 6365 5284 6377 5287
rect 4948 5256 6377 5284
rect 4948 5244 4954 5256
rect 6365 5253 6377 5256
rect 6411 5253 6423 5287
rect 6546 5284 6552 5296
rect 6507 5256 6552 5284
rect 6365 5247 6423 5253
rect 6546 5244 6552 5256
rect 6604 5244 6610 5296
rect 6730 5244 6736 5296
rect 6788 5284 6794 5296
rect 8570 5284 8576 5296
rect 6788 5256 8576 5284
rect 6788 5244 6794 5256
rect 8570 5244 8576 5256
rect 8628 5244 8634 5296
rect 9214 5284 9220 5296
rect 9175 5256 9220 5284
rect 9214 5244 9220 5256
rect 9272 5244 9278 5296
rect 13630 5244 13636 5296
rect 13688 5284 13694 5296
rect 17126 5284 17132 5296
rect 13688 5256 17132 5284
rect 13688 5244 13694 5256
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 5258 5216 5264 5228
rect 4203 5188 5264 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 5169 5151 5227 5157
rect 5169 5148 5181 5151
rect 4304 5120 5181 5148
rect 4304 5108 4310 5120
rect 5169 5117 5181 5120
rect 5215 5117 5227 5151
rect 5276 5148 5304 5176
rect 6822 5148 6828 5160
rect 5276 5120 6828 5148
rect 5169 5111 5227 5117
rect 6822 5108 6828 5120
rect 6880 5148 6886 5160
rect 7208 5148 7236 5179
rect 8202 5176 8208 5228
rect 8260 5216 8266 5228
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 8260 5188 9137 5216
rect 8260 5176 8266 5188
rect 9125 5185 9137 5188
rect 9171 5216 9183 5219
rect 9766 5216 9772 5228
rect 9171 5188 9772 5216
rect 9171 5185 9183 5188
rect 9125 5179 9183 5185
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 6880 5120 7236 5148
rect 6880 5108 6886 5120
rect 6638 4972 6644 5024
rect 6696 5012 6702 5024
rect 6733 5015 6791 5021
rect 6733 5012 6745 5015
rect 6696 4984 6745 5012
rect 6696 4972 6702 4984
rect 6733 4981 6745 4984
rect 6779 4981 6791 5015
rect 6733 4975 6791 4981
rect 3036 4922 9844 4944
rect 3036 4870 7566 4922
rect 7618 4870 7630 4922
rect 7682 4870 7694 4922
rect 7746 4870 7758 4922
rect 7810 4870 7822 4922
rect 7874 4870 9844 4922
rect 3036 4848 9844 4870
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 3970 4808 3976 4820
rect 3651 4780 3976 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 4706 4808 4712 4820
rect 4667 4780 4712 4808
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5350 4808 5356 4820
rect 5307 4780 5356 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 6733 4811 6791 4817
rect 6733 4808 6745 4811
rect 6144 4780 6745 4808
rect 6144 4768 6150 4780
rect 6733 4777 6745 4780
rect 6779 4777 6791 4811
rect 7374 4808 7380 4820
rect 7335 4780 7380 4808
rect 6733 4771 6791 4777
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 8352 4780 8401 4808
rect 8352 4768 8358 4780
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 8389 4771 8447 4777
rect 9217 4811 9275 4817
rect 9217 4777 9229 4811
rect 9263 4808 9275 4811
rect 9398 4808 9404 4820
rect 9263 4780 9404 4808
rect 9263 4777 9275 4780
rect 9217 4771 9275 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 17402 4808 17408 4820
rect 12400 4780 17408 4808
rect 12400 4768 12406 4780
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 474 4700 480 4752
rect 532 4740 538 4752
rect 5534 4740 5540 4752
rect 532 4712 5540 4740
rect 532 4700 538 4712
rect 5534 4700 5540 4712
rect 5592 4700 5598 4752
rect 2038 4632 2044 4684
rect 2096 4672 2102 4684
rect 2590 4672 2596 4684
rect 2096 4644 2596 4672
rect 2096 4632 2102 4644
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 8110 4672 8116 4684
rect 7300 4644 8116 4672
rect 1210 4564 1216 4616
rect 1268 4604 1274 4616
rect 2866 4604 2872 4616
rect 1268 4576 2872 4604
rect 1268 4564 1274 4576
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 3510 4604 3516 4616
rect 3471 4576 3516 4604
rect 3510 4564 3516 4576
rect 3568 4564 3574 4616
rect 4522 4604 4528 4616
rect 4483 4576 4528 4604
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 5169 4607 5227 4613
rect 5169 4604 5181 4607
rect 4948 4576 5181 4604
rect 4948 4564 4954 4576
rect 5169 4573 5181 4576
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 5442 4604 5448 4616
rect 5399 4576 5448 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 6178 4604 6184 4616
rect 6139 4576 6184 4604
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 6822 4604 6828 4616
rect 6783 4576 6828 4604
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 7300 4613 7328 4644
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 7432 4576 7481 4604
rect 7432 4564 7438 4576
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 8570 4604 8576 4616
rect 8531 4576 8576 4604
rect 7469 4567 7527 4573
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4604 9091 4607
rect 9674 4604 9680 4616
rect 9079 4576 9680 4604
rect 9079 4573 9091 4576
rect 9033 4567 9091 4573
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 842 4496 848 4548
rect 900 4536 906 4548
rect 2958 4536 2964 4548
rect 900 4508 2964 4536
rect 900 4496 906 4508
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4468 6055 4471
rect 6730 4468 6736 4480
rect 6043 4440 6736 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 3036 4378 9844 4400
rect 3036 4326 3566 4378
rect 3618 4326 3630 4378
rect 3682 4326 3694 4378
rect 3746 4326 3758 4378
rect 3810 4326 3822 4378
rect 3874 4326 8566 4378
rect 8618 4326 8630 4378
rect 8682 4326 8694 4378
rect 8746 4326 8758 4378
rect 8810 4326 8822 4378
rect 8874 4326 9844 4378
rect 3036 4304 9844 4326
rect 3510 4224 3516 4276
rect 3568 4264 3574 4276
rect 5718 4264 5724 4276
rect 3568 4236 5724 4264
rect 3568 4224 3574 4236
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 7009 4267 7067 4273
rect 7009 4233 7021 4267
rect 7055 4264 7067 4267
rect 7098 4264 7104 4276
rect 7055 4236 7104 4264
rect 7055 4233 7067 4236
rect 7009 4227 7067 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 7374 4224 7380 4276
rect 7432 4264 7438 4276
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 7432 4236 7573 4264
rect 7432 4224 7438 4236
rect 7561 4233 7573 4236
rect 7607 4233 7619 4267
rect 7561 4227 7619 4233
rect 10870 4224 10876 4276
rect 10928 4264 10934 4276
rect 18230 4264 18236 4276
rect 10928 4236 18236 4264
rect 10928 4224 10934 4236
rect 18230 4224 18236 4236
rect 18288 4224 18294 4276
rect 3418 4156 3424 4208
rect 3476 4196 3482 4208
rect 3476 4168 4108 4196
rect 3476 4156 3482 4168
rect 2682 4088 2688 4140
rect 2740 4128 2746 4140
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 2740 4100 3709 4128
rect 2740 4088 2746 4100
rect 3697 4097 3709 4100
rect 3743 4097 3755 4131
rect 4080 4128 4108 4168
rect 6454 4156 6460 4208
rect 6512 4196 6518 4208
rect 7392 4196 7420 4224
rect 6512 4168 6960 4196
rect 6512 4156 6518 4168
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 4080 4100 4813 4128
rect 3697 4091 3755 4097
rect 4801 4097 4813 4100
rect 4847 4128 4859 4131
rect 4890 4128 4896 4140
rect 4847 4100 4896 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 5629 4131 5687 4137
rect 5629 4128 5641 4131
rect 5592 4100 5641 4128
rect 5592 4088 5598 4100
rect 5629 4097 5641 4100
rect 5675 4097 5687 4131
rect 6086 4128 6092 4140
rect 6047 4100 6092 4128
rect 5629 4091 5687 4097
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 6270 4128 6276 4140
rect 6231 4100 6276 4128
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 6546 4088 6552 4140
rect 6604 4128 6610 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6604 4100 6837 4128
rect 6604 4088 6610 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 4062 4060 4068 4072
rect 4023 4032 4068 4060
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 6181 4063 6239 4069
rect 6181 4060 6193 4063
rect 5868 4032 6193 4060
rect 5868 4020 5874 4032
rect 6181 4029 6193 4032
rect 6227 4029 6239 4063
rect 6932 4060 6960 4168
rect 7024 4168 7420 4196
rect 7024 4137 7052 4168
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7668 4060 7696 4091
rect 8478 4088 8484 4140
rect 8536 4128 8542 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8536 4100 9045 4128
rect 8536 4088 8542 4100
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 6932 4032 7696 4060
rect 6181 4023 6239 4029
rect 4893 3995 4951 4001
rect 4893 3961 4905 3995
rect 4939 3992 4951 3995
rect 4982 3992 4988 4004
rect 4939 3964 4988 3992
rect 4939 3961 4951 3964
rect 4893 3955 4951 3961
rect 4982 3952 4988 3964
rect 5040 3952 5046 4004
rect 6270 3952 6276 4004
rect 6328 3992 6334 4004
rect 10778 3992 10784 4004
rect 6328 3964 10784 3992
rect 6328 3952 6334 3964
rect 10778 3952 10784 3964
rect 10836 3952 10842 4004
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4706 3924 4712 3936
rect 4120 3896 4712 3924
rect 4120 3884 4126 3896
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 5442 3924 5448 3936
rect 5403 3896 5448 3924
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 9214 3924 9220 3936
rect 9175 3896 9220 3924
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 16850 3924 16856 3936
rect 13872 3896 16856 3924
rect 13872 3884 13878 3896
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 3036 3834 9844 3856
rect 3036 3782 7566 3834
rect 7618 3782 7630 3834
rect 7682 3782 7694 3834
rect 7746 3782 7758 3834
rect 7810 3782 7822 3834
rect 7874 3782 9844 3834
rect 3036 3760 9844 3782
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 3605 3723 3663 3729
rect 3605 3720 3617 3723
rect 3108 3692 3617 3720
rect 3108 3680 3114 3692
rect 3605 3689 3617 3692
rect 3651 3689 3663 3723
rect 3605 3683 3663 3689
rect 4341 3723 4399 3729
rect 4341 3689 4353 3723
rect 4387 3720 4399 3723
rect 4614 3720 4620 3732
rect 4387 3692 4620 3720
rect 4387 3689 4399 3692
rect 4341 3683 4399 3689
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 4985 3723 5043 3729
rect 4985 3689 4997 3723
rect 5031 3720 5043 3723
rect 5074 3720 5080 3732
rect 5031 3692 5080 3720
rect 5031 3689 5043 3692
rect 4985 3683 5043 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 5994 3720 6000 3732
rect 5955 3692 6000 3720
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 4706 3584 4712 3596
rect 3712 3556 4712 3584
rect 2958 3476 2964 3528
rect 3016 3516 3022 3528
rect 3712 3525 3740 3556
rect 4706 3544 4712 3556
rect 4764 3584 4770 3596
rect 6178 3584 6184 3596
rect 4764 3556 6184 3584
rect 4764 3544 4770 3556
rect 6178 3544 6184 3556
rect 6236 3584 6242 3596
rect 6236 3556 7236 3584
rect 6236 3544 6242 3556
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 3016 3488 3525 3516
rect 3016 3476 3022 3488
rect 3513 3485 3525 3488
rect 3559 3485 3571 3519
rect 3513 3479 3571 3485
rect 3697 3519 3755 3525
rect 3697 3485 3709 3519
rect 3743 3485 3755 3519
rect 4154 3516 4160 3528
rect 4115 3488 4160 3516
rect 3697 3479 3755 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4890 3516 4896 3528
rect 4851 3488 4896 3516
rect 4890 3476 4896 3488
rect 4948 3516 4954 3528
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 4948 3488 6101 3516
rect 4948 3476 4954 3488
rect 6089 3485 6101 3488
rect 6135 3516 6147 3519
rect 6914 3516 6920 3528
rect 6135 3488 6920 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 7208 3525 7236 3556
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 9950 3584 9956 3596
rect 8352 3556 9956 3584
rect 8352 3544 8358 3556
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 7193 3519 7251 3525
rect 7064 3488 7109 3516
rect 7064 3476 7070 3488
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 8202 3516 8208 3528
rect 8163 3488 8208 3516
rect 7193 3479 7251 3485
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 9033 3519 9091 3525
rect 9033 3516 9045 3519
rect 8996 3488 9045 3516
rect 8996 3476 9002 3488
rect 9033 3485 9045 3488
rect 9079 3485 9091 3519
rect 9033 3479 9091 3485
rect 7926 3408 7932 3460
rect 7984 3448 7990 3460
rect 11790 3448 11796 3460
rect 7984 3420 11796 3448
rect 7984 3408 7990 3420
rect 11790 3408 11796 3420
rect 11848 3408 11854 3460
rect 12250 3408 12256 3460
rect 12308 3448 12314 3460
rect 12894 3448 12900 3460
rect 12308 3420 12900 3448
rect 12308 3408 12314 3420
rect 12894 3408 12900 3420
rect 12952 3408 12958 3460
rect 7190 3380 7196 3392
rect 7151 3352 7196 3380
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 8168 3352 8309 3380
rect 8168 3340 8174 3352
rect 8297 3349 8309 3352
rect 8343 3349 8355 3383
rect 9214 3380 9220 3392
rect 9175 3352 9220 3380
rect 8297 3343 8355 3349
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 3036 3290 9844 3312
rect 3036 3238 3566 3290
rect 3618 3238 3630 3290
rect 3682 3238 3694 3290
rect 3746 3238 3758 3290
rect 3810 3238 3822 3290
rect 3874 3238 8566 3290
rect 8618 3238 8630 3290
rect 8682 3238 8694 3290
rect 8746 3238 8758 3290
rect 8810 3238 8822 3290
rect 8874 3238 9844 3290
rect 3036 3216 9844 3238
rect 4801 3179 4859 3185
rect 4801 3145 4813 3179
rect 4847 3176 4859 3179
rect 5258 3176 5264 3188
rect 4847 3148 5264 3176
rect 4847 3145 4859 3148
rect 4801 3139 4859 3145
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 6181 3179 6239 3185
rect 6181 3145 6193 3179
rect 6227 3176 6239 3179
rect 6270 3176 6276 3188
rect 6227 3148 6276 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 7466 3176 7472 3188
rect 7239 3148 7472 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 8018 3176 8024 3188
rect 7883 3148 8024 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 9858 3176 9864 3188
rect 8220 3148 9864 3176
rect 3970 3108 3976 3120
rect 3931 3080 3976 3108
rect 3970 3068 3976 3080
rect 4028 3068 4034 3120
rect 6638 3068 6644 3120
rect 6696 3108 6702 3120
rect 6696 3080 7696 3108
rect 6696 3068 6702 3080
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 2924 3012 3617 3040
rect 2924 3000 2930 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 4706 3040 4712 3052
rect 3752 3012 4712 3040
rect 3752 3000 3758 3012
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3040 4951 3043
rect 5166 3040 5172 3052
rect 4939 3012 5172 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5350 3040 5356 3052
rect 5311 3012 5356 3040
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3040 6055 3043
rect 6362 3040 6368 3052
rect 6043 3012 6368 3040
rect 6043 3009 6055 3012
rect 5997 3003 6055 3009
rect 5552 2972 5580 3003
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 7668 3049 7696 3080
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3009 7711 3043
rect 7653 3003 7711 3009
rect 6546 2972 6552 2984
rect 5552 2944 6552 2972
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 7024 2972 7052 3003
rect 8220 2972 8248 3148
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 10042 3108 10048 3120
rect 8680 3080 10048 3108
rect 8680 3049 8708 3080
rect 10042 3068 10048 3080
rect 10100 3068 10106 3120
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 7024 2944 8248 2972
rect 7834 2864 7840 2916
rect 7892 2904 7898 2916
rect 8496 2904 8524 3003
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 9125 3043 9183 3049
rect 9125 3040 9137 3043
rect 9088 3012 9137 3040
rect 9088 3000 9094 3012
rect 9125 3009 9137 3012
rect 9171 3009 9183 3043
rect 9125 3003 9183 3009
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 8570 2932 8576 2984
rect 8628 2972 8634 2984
rect 9324 2972 9352 3003
rect 8628 2944 9352 2972
rect 8628 2932 8634 2944
rect 9214 2904 9220 2916
rect 7892 2876 8524 2904
rect 9175 2876 9220 2904
rect 7892 2864 7898 2876
rect 9214 2864 9220 2876
rect 9272 2864 9278 2916
rect 5445 2839 5503 2845
rect 5445 2805 5457 2839
rect 5491 2836 5503 2839
rect 5534 2836 5540 2848
rect 5491 2808 5540 2836
rect 5491 2805 5503 2808
rect 5445 2799 5503 2805
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 8202 2796 8208 2848
rect 8260 2836 8266 2848
rect 8573 2839 8631 2845
rect 8573 2836 8585 2839
rect 8260 2808 8585 2836
rect 8260 2796 8266 2808
rect 8573 2805 8585 2808
rect 8619 2805 8631 2839
rect 8573 2799 8631 2805
rect 3036 2746 9844 2768
rect 3036 2694 7566 2746
rect 7618 2694 7630 2746
rect 7682 2694 7694 2746
rect 7746 2694 7758 2746
rect 7810 2694 7822 2746
rect 7874 2694 9844 2746
rect 17586 2728 17592 2780
rect 17644 2768 17650 2780
rect 17954 2768 17960 2780
rect 17644 2740 17960 2768
rect 17644 2728 17650 2740
rect 17954 2728 17960 2740
rect 18012 2728 18018 2780
rect 3036 2672 9844 2694
rect 3605 2635 3663 2641
rect 3605 2601 3617 2635
rect 3651 2632 3663 2635
rect 3970 2632 3976 2644
rect 3651 2604 3976 2632
rect 3651 2601 3663 2604
rect 3605 2595 3663 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 8570 2632 8576 2644
rect 8531 2604 8576 2632
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 9398 2632 9404 2644
rect 9171 2604 9404 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 5626 2524 5632 2576
rect 5684 2564 5690 2576
rect 5684 2536 6776 2564
rect 5684 2524 5690 2536
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 5592 2468 6592 2496
rect 5592 2456 5598 2468
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 2832 2400 3525 2428
rect 2832 2388 2838 2400
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3694 2428 3700 2440
rect 3655 2400 3700 2428
rect 3513 2391 3571 2397
rect 3694 2388 3700 2400
rect 3752 2388 3758 2440
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 5902 2428 5908 2440
rect 5863 2400 5908 2428
rect 4893 2391 4951 2397
rect 4908 2360 4936 2391
rect 5902 2388 5908 2400
rect 5960 2388 5966 2440
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2428 6147 2431
rect 6270 2428 6276 2440
rect 6135 2400 6276 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 6564 2437 6592 2468
rect 6748 2437 6776 2536
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2397 6791 2431
rect 7190 2428 7196 2440
rect 7151 2400 7196 2428
rect 6733 2391 6791 2397
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2428 7435 2431
rect 8202 2428 8208 2440
rect 7423 2400 8208 2428
rect 7423 2397 7435 2400
rect 7377 2391 7435 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2428 8723 2431
rect 9122 2428 9128 2440
rect 8711 2400 9128 2428
rect 8711 2397 8723 2400
rect 8665 2391 8723 2397
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 9306 2428 9312 2440
rect 9267 2400 9312 2428
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 8294 2360 8300 2372
rect 4908 2332 8300 2360
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 4706 2292 4712 2304
rect 4667 2264 4712 2292
rect 4706 2252 4712 2264
rect 4764 2252 4770 2304
rect 5994 2292 6000 2304
rect 5955 2264 6000 2292
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 6730 2292 6736 2304
rect 6691 2264 6736 2292
rect 6730 2252 6736 2264
rect 6788 2252 6794 2304
rect 6822 2252 6828 2304
rect 6880 2292 6886 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 6880 2264 7297 2292
rect 6880 2252 6886 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 3036 2202 9844 2224
rect 3036 2150 3566 2202
rect 3618 2150 3630 2202
rect 3682 2150 3694 2202
rect 3746 2150 3758 2202
rect 3810 2150 3822 2202
rect 3874 2150 8566 2202
rect 8618 2150 8630 2202
rect 8682 2150 8694 2202
rect 8746 2150 8758 2202
rect 8810 2150 8822 2202
rect 8874 2150 9844 2202
rect 3036 2128 9844 2150
rect 3697 2091 3755 2097
rect 3697 2057 3709 2091
rect 3743 2088 3755 2091
rect 4062 2088 4068 2100
rect 3743 2060 4068 2088
rect 3743 2057 3755 2060
rect 3697 2051 3755 2057
rect 4062 2048 4068 2060
rect 4120 2048 4126 2100
rect 4338 2088 4344 2100
rect 4299 2060 4344 2088
rect 4338 2048 4344 2060
rect 4396 2048 4402 2100
rect 4985 2091 5043 2097
rect 4985 2057 4997 2091
rect 5031 2088 5043 2091
rect 5350 2088 5356 2100
rect 5031 2060 5356 2088
rect 5031 2057 5043 2060
rect 4985 2051 5043 2057
rect 5350 2048 5356 2060
rect 5408 2048 5414 2100
rect 5626 2088 5632 2100
rect 5587 2060 5632 2088
rect 5626 2048 5632 2060
rect 5684 2048 5690 2100
rect 6638 2048 6644 2100
rect 6696 2088 6702 2100
rect 6733 2091 6791 2097
rect 6733 2088 6745 2091
rect 6696 2060 6745 2088
rect 6696 2048 6702 2060
rect 6733 2057 6745 2060
rect 6779 2057 6791 2091
rect 6733 2051 6791 2057
rect 8665 2091 8723 2097
rect 8665 2057 8677 2091
rect 8711 2088 8723 2091
rect 8938 2088 8944 2100
rect 8711 2060 8944 2088
rect 8711 2057 8723 2060
rect 8665 2051 8723 2057
rect 8938 2048 8944 2060
rect 8996 2048 9002 2100
rect 9214 2088 9220 2100
rect 9175 2060 9220 2088
rect 9214 2048 9220 2060
rect 9272 2048 9278 2100
rect 8110 2020 8116 2032
rect 6932 1992 8116 2020
rect 3418 1912 3424 1964
rect 3476 1952 3482 1964
rect 3513 1955 3571 1961
rect 3513 1952 3525 1955
rect 3476 1924 3525 1952
rect 3476 1912 3482 1924
rect 3513 1921 3525 1924
rect 3559 1921 3571 1955
rect 4154 1952 4160 1964
rect 4115 1924 4160 1952
rect 3513 1915 3571 1921
rect 4154 1912 4160 1924
rect 4212 1912 4218 1964
rect 4798 1952 4804 1964
rect 4759 1924 4804 1952
rect 4798 1912 4804 1924
rect 4856 1912 4862 1964
rect 4985 1955 5043 1961
rect 4985 1921 4997 1955
rect 5031 1921 5043 1955
rect 5442 1952 5448 1964
rect 5403 1924 5448 1952
rect 4985 1915 5043 1921
rect 5000 1884 5028 1915
rect 5442 1912 5448 1924
rect 5500 1912 5506 1964
rect 6086 1952 6092 1964
rect 6047 1924 6092 1952
rect 6086 1912 6092 1924
rect 6144 1912 6150 1964
rect 6270 1952 6276 1964
rect 6231 1924 6276 1952
rect 6270 1912 6276 1924
rect 6328 1912 6334 1964
rect 6733 1955 6791 1961
rect 6733 1921 6745 1955
rect 6779 1952 6791 1955
rect 6822 1952 6828 1964
rect 6779 1924 6828 1952
rect 6779 1921 6791 1924
rect 6733 1915 6791 1921
rect 6822 1912 6828 1924
rect 6880 1912 6886 1964
rect 6932 1961 6960 1992
rect 8110 1980 8116 1992
rect 8168 1980 8174 2032
rect 6917 1955 6975 1961
rect 6917 1921 6929 1955
rect 6963 1921 6975 1955
rect 6917 1915 6975 1921
rect 7006 1912 7012 1964
rect 7064 1952 7070 1964
rect 7377 1955 7435 1961
rect 7377 1952 7389 1955
rect 7064 1924 7389 1952
rect 7064 1912 7070 1924
rect 7377 1921 7389 1924
rect 7423 1921 7435 1955
rect 7377 1915 7435 1921
rect 8481 1955 8539 1961
rect 8481 1921 8493 1955
rect 8527 1952 8539 1955
rect 9030 1952 9036 1964
rect 8527 1924 9036 1952
rect 8527 1921 8539 1924
rect 8481 1915 8539 1921
rect 9030 1912 9036 1924
rect 9088 1912 9094 1964
rect 9306 1952 9312 1964
rect 9267 1924 9312 1952
rect 9306 1912 9312 1924
rect 9364 1912 9370 1964
rect 6288 1884 6316 1912
rect 5000 1856 6316 1884
rect 7466 1816 7472 1828
rect 7427 1788 7472 1816
rect 7466 1776 7472 1788
rect 7524 1776 7530 1828
rect 6178 1748 6184 1760
rect 6139 1720 6184 1748
rect 6178 1708 6184 1720
rect 6236 1708 6242 1760
rect 3036 1658 9844 1680
rect 3036 1606 7566 1658
rect 7618 1606 7630 1658
rect 7682 1606 7694 1658
rect 7746 1606 7758 1658
rect 7810 1606 7822 1658
rect 7874 1606 9844 1658
rect 3036 1584 9844 1606
rect 750 1504 756 1556
rect 808 1544 814 1556
rect 4798 1544 4804 1556
rect 808 1516 4804 1544
rect 808 1504 814 1516
rect 4798 1504 4804 1516
rect 4856 1504 4862 1556
rect 6546 1504 6552 1556
rect 6604 1544 6610 1556
rect 6641 1547 6699 1553
rect 6641 1544 6653 1547
rect 6604 1516 6653 1544
rect 6604 1504 6610 1516
rect 6641 1513 6653 1516
rect 6687 1513 6699 1547
rect 6641 1507 6699 1513
rect 4522 1368 4528 1420
rect 4580 1408 4586 1420
rect 4580 1380 5212 1408
rect 4580 1368 4586 1380
rect 3602 1340 3608 1352
rect 3563 1312 3608 1340
rect 3602 1300 3608 1312
rect 3660 1300 3666 1352
rect 3697 1343 3755 1349
rect 3697 1309 3709 1343
rect 3743 1309 3755 1343
rect 4154 1340 4160 1352
rect 4115 1312 4160 1340
rect 3697 1303 3755 1309
rect 3234 1232 3240 1284
rect 3292 1272 3298 1284
rect 3712 1272 3740 1303
rect 4154 1300 4160 1312
rect 4212 1300 4218 1352
rect 4801 1343 4859 1349
rect 4801 1309 4813 1343
rect 4847 1340 4859 1343
rect 5074 1340 5080 1352
rect 4847 1312 5080 1340
rect 4847 1309 4859 1312
rect 4801 1303 4859 1309
rect 5074 1300 5080 1312
rect 5132 1300 5138 1352
rect 5184 1340 5212 1380
rect 5905 1343 5963 1349
rect 5905 1340 5917 1343
rect 5184 1312 5917 1340
rect 5905 1309 5917 1312
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 6089 1343 6147 1349
rect 6089 1309 6101 1343
rect 6135 1340 6147 1343
rect 6270 1340 6276 1352
rect 6135 1312 6276 1340
rect 6135 1309 6147 1312
rect 6089 1303 6147 1309
rect 6270 1300 6276 1312
rect 6328 1300 6334 1352
rect 6730 1340 6736 1352
rect 6691 1312 6736 1340
rect 6730 1300 6736 1312
rect 6788 1300 6794 1352
rect 7374 1340 7380 1352
rect 7335 1312 7380 1340
rect 7374 1300 7380 1312
rect 7432 1300 7438 1352
rect 4062 1272 4068 1284
rect 3292 1244 4068 1272
rect 3292 1232 3298 1244
rect 4062 1232 4068 1244
rect 4120 1232 4126 1284
rect 7285 1275 7343 1281
rect 7285 1241 7297 1275
rect 7331 1272 7343 1275
rect 8202 1272 8208 1284
rect 7331 1244 8208 1272
rect 7331 1241 7343 1244
rect 7285 1235 7343 1241
rect 8202 1232 8208 1244
rect 8260 1232 8266 1284
rect 4338 1204 4344 1216
rect 4299 1176 4344 1204
rect 4338 1164 4344 1176
rect 4396 1164 4402 1216
rect 4890 1204 4896 1216
rect 4851 1176 4896 1204
rect 4890 1164 4896 1176
rect 4948 1164 4954 1216
rect 5994 1204 6000 1216
rect 5955 1176 6000 1204
rect 5994 1164 6000 1176
rect 6052 1164 6058 1216
rect 3036 1114 9844 1136
rect 3036 1062 3566 1114
rect 3618 1062 3630 1114
rect 3682 1062 3694 1114
rect 3746 1062 3758 1114
rect 3810 1062 3822 1114
rect 3874 1062 8566 1114
rect 8618 1062 8630 1114
rect 8682 1062 8694 1114
rect 8746 1062 8758 1114
rect 8810 1062 8822 1114
rect 8874 1062 9844 1114
rect 3036 1040 9844 1062
<< via1 >>
rect 13636 16668 13688 16720
rect 15292 16668 15344 16720
rect 2566 15750 2618 15802
rect 2630 15750 2682 15802
rect 2694 15750 2746 15802
rect 2758 15750 2810 15802
rect 2822 15750 2874 15802
rect 7566 15750 7618 15802
rect 7630 15750 7682 15802
rect 7694 15750 7746 15802
rect 7758 15750 7810 15802
rect 7822 15750 7874 15802
rect 2412 15648 2464 15700
rect 5724 15691 5776 15700
rect 5724 15657 5733 15691
rect 5733 15657 5767 15691
rect 5767 15657 5776 15691
rect 5724 15648 5776 15657
rect 4712 15555 4764 15564
rect 4712 15521 4721 15555
rect 4721 15521 4755 15555
rect 4755 15521 4764 15555
rect 4712 15512 4764 15521
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 1124 15376 1176 15428
rect 3056 15444 3108 15496
rect 4068 15444 4120 15496
rect 5448 15444 5500 15496
rect 6184 15444 6236 15496
rect 8392 15487 8444 15496
rect 8392 15453 8401 15487
rect 8401 15453 8435 15487
rect 8435 15453 8444 15487
rect 8392 15444 8444 15453
rect 9036 15444 9088 15496
rect 3148 15419 3200 15428
rect 3148 15385 3157 15419
rect 3157 15385 3191 15419
rect 3191 15385 3200 15419
rect 3148 15376 3200 15385
rect 7840 15376 7892 15428
rect 8116 15419 8168 15428
rect 8116 15385 8125 15419
rect 8125 15385 8159 15419
rect 8159 15385 8168 15419
rect 8116 15376 8168 15385
rect 1308 15308 1360 15360
rect 2780 15308 2832 15360
rect 5356 15308 5408 15360
rect 9128 15351 9180 15360
rect 9128 15317 9137 15351
rect 9137 15317 9171 15351
rect 9171 15317 9180 15351
rect 9128 15308 9180 15317
rect 3566 15206 3618 15258
rect 3630 15206 3682 15258
rect 3694 15206 3746 15258
rect 3758 15206 3810 15258
rect 3822 15206 3874 15258
rect 8566 15206 8618 15258
rect 8630 15206 8682 15258
rect 8694 15206 8746 15258
rect 8758 15206 8810 15258
rect 8822 15206 8874 15258
rect 13636 15240 13688 15292
rect 16488 15240 16540 15292
rect 1676 15104 1728 15156
rect 940 15036 992 15088
rect 5540 15104 5592 15156
rect 17914 15104 17966 15156
rect 18788 15104 18840 15156
rect 1584 14968 1636 15020
rect 1676 15011 1728 15020
rect 1676 14977 1685 15011
rect 1685 14977 1719 15011
rect 1719 14977 1728 15011
rect 1676 14968 1728 14977
rect 2320 14968 2372 15020
rect 7840 15036 7892 15088
rect 8208 15036 8260 15088
rect 1400 14900 1452 14952
rect 3516 14968 3568 15020
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 8944 15011 8996 15020
rect 8944 14977 8953 15011
rect 8953 14977 8987 15011
rect 8987 14977 8996 15011
rect 8944 14968 8996 14977
rect 5724 14943 5776 14952
rect 5724 14909 5733 14943
rect 5733 14909 5767 14943
rect 5767 14909 5776 14943
rect 5724 14900 5776 14909
rect 8392 14943 8444 14952
rect 8392 14909 8401 14943
rect 8401 14909 8435 14943
rect 8435 14909 8444 14943
rect 8392 14900 8444 14909
rect 2780 14875 2832 14884
rect 2780 14841 2789 14875
rect 2789 14841 2823 14875
rect 2823 14841 2832 14875
rect 2780 14832 2832 14841
rect 4160 14832 4212 14884
rect 13636 14832 13688 14884
rect 17408 14832 17460 14884
rect 296 14764 348 14816
rect 4068 14764 4120 14816
rect 4528 14764 4580 14816
rect 9128 14807 9180 14816
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 13820 14764 13872 14816
rect 15292 14764 15344 14816
rect 2566 14662 2618 14714
rect 2630 14662 2682 14714
rect 2694 14662 2746 14714
rect 2758 14662 2810 14714
rect 2822 14662 2874 14714
rect 7566 14662 7618 14714
rect 7630 14662 7682 14714
rect 7694 14662 7746 14714
rect 7758 14662 7810 14714
rect 7822 14662 7874 14714
rect 13636 14696 13688 14748
rect 14188 14696 14240 14748
rect 13636 14560 13688 14612
rect 14832 14560 14884 14612
rect 3976 14492 4028 14544
rect 4436 14535 4488 14544
rect 4436 14501 4445 14535
rect 4445 14501 4479 14535
rect 4479 14501 4488 14535
rect 4436 14492 4488 14501
rect 5264 14467 5316 14476
rect 5264 14433 5273 14467
rect 5273 14433 5307 14467
rect 5307 14433 5316 14467
rect 5264 14424 5316 14433
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3976 14399 4028 14408
rect 3240 14356 3292 14365
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 4712 14356 4764 14408
rect 6460 14356 6512 14408
rect 8208 14356 8260 14408
rect 8392 14424 8444 14476
rect 15384 14424 15436 14476
rect 9220 14356 9272 14408
rect 15200 14356 15252 14408
rect 17592 14356 17644 14408
rect 2504 14288 2556 14340
rect 3516 14288 3568 14340
rect 5356 14288 5408 14340
rect 7380 14288 7432 14340
rect 9404 14288 9456 14340
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 3976 14220 4028 14272
rect 8484 14220 8536 14272
rect 9312 14263 9364 14272
rect 9312 14229 9321 14263
rect 9321 14229 9355 14263
rect 9355 14229 9364 14263
rect 9312 14220 9364 14229
rect 3566 14118 3618 14170
rect 3630 14118 3682 14170
rect 3694 14118 3746 14170
rect 3758 14118 3810 14170
rect 3822 14118 3874 14170
rect 8566 14118 8618 14170
rect 8630 14118 8682 14170
rect 8694 14118 8746 14170
rect 8758 14118 8810 14170
rect 8822 14118 8874 14170
rect 12808 14152 12860 14204
rect 17132 14152 17184 14204
rect 5448 14059 5500 14068
rect 5448 14025 5457 14059
rect 5457 14025 5491 14059
rect 5491 14025 5500 14059
rect 5448 14016 5500 14025
rect 4068 13948 4120 14000
rect 5080 13948 5132 14000
rect 1492 13880 1544 13932
rect 2412 13880 2464 13932
rect 2780 13880 2832 13932
rect 4528 13923 4580 13932
rect 4528 13889 4537 13923
rect 4537 13889 4571 13923
rect 4571 13889 4580 13923
rect 4528 13880 4580 13889
rect 4896 13923 4948 13932
rect 4896 13889 4905 13923
rect 4905 13889 4939 13923
rect 4939 13889 4948 13923
rect 4896 13880 4948 13889
rect 5448 13880 5500 13932
rect 2964 13744 3016 13796
rect 9128 14016 9180 14068
rect 8116 13948 8168 14000
rect 8484 13880 8536 13932
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 6644 13812 6696 13821
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 8944 13812 8996 13821
rect 6000 13744 6052 13796
rect 1768 13676 1820 13728
rect 2504 13676 2556 13728
rect 3056 13676 3108 13728
rect 8024 13676 8076 13728
rect 2566 13574 2618 13626
rect 2630 13574 2682 13626
rect 2694 13574 2746 13626
rect 2758 13574 2810 13626
rect 2822 13574 2874 13626
rect 7566 13574 7618 13626
rect 7630 13574 7682 13626
rect 7694 13574 7746 13626
rect 7758 13574 7810 13626
rect 7822 13574 7874 13626
rect 13728 13540 13780 13592
rect 16028 13540 16080 13592
rect 17914 13540 17966 13592
rect 18972 13540 19024 13592
rect 13820 13472 13872 13524
rect 18328 13472 18380 13524
rect 15752 13404 15804 13456
rect 112 13336 164 13388
rect 1400 13336 1452 13388
rect 5448 13336 5500 13388
rect 3056 13268 3108 13320
rect 4068 13268 4120 13320
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 7012 13268 7064 13277
rect 8392 13268 8444 13320
rect 1400 13200 1452 13252
rect 6644 13200 6696 13252
rect 1584 13132 1636 13184
rect 15476 13200 15528 13252
rect 3566 13030 3618 13082
rect 3630 13030 3682 13082
rect 3694 13030 3746 13082
rect 3758 13030 3810 13082
rect 3822 13030 3874 13082
rect 8566 13030 8618 13082
rect 8630 13030 8682 13082
rect 8694 13030 8746 13082
rect 8758 13030 8810 13082
rect 8822 13030 8874 13082
rect 8300 12971 8352 12980
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 13820 12928 13872 12980
rect 17316 12928 17368 12980
rect 3516 12860 3568 12912
rect 1768 12792 1820 12844
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 4436 12835 4488 12844
rect 4436 12801 4445 12835
rect 4445 12801 4479 12835
rect 4479 12801 4488 12835
rect 4436 12792 4488 12801
rect 5264 12792 5316 12844
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 7932 12792 7984 12844
rect 15016 12792 15068 12844
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 5816 12724 5868 12776
rect 7196 12724 7248 12776
rect 13452 12656 13504 12708
rect 15200 12656 15252 12708
rect 848 12588 900 12640
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 7932 12588 7984 12640
rect 9496 12588 9548 12640
rect 2566 12486 2618 12538
rect 2630 12486 2682 12538
rect 2694 12486 2746 12538
rect 2758 12486 2810 12538
rect 2822 12486 2874 12538
rect 7566 12486 7618 12538
rect 7630 12486 7682 12538
rect 7694 12486 7746 12538
rect 7758 12486 7810 12538
rect 7822 12486 7874 12538
rect 13820 12520 13872 12572
rect 15936 12520 15988 12572
rect 664 12384 716 12436
rect 1216 12384 1268 12436
rect 2412 12248 2464 12300
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 3424 12180 3476 12232
rect 3056 12112 3108 12164
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 2964 12044 3016 12096
rect 4068 12180 4120 12232
rect 4252 12180 4304 12232
rect 4712 12180 4764 12232
rect 6276 12223 6328 12232
rect 6276 12189 6285 12223
rect 6285 12189 6319 12223
rect 6319 12189 6328 12223
rect 6276 12180 6328 12189
rect 7196 12180 7248 12232
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 8760 12180 8812 12232
rect 12348 12180 12400 12232
rect 12992 12180 13044 12232
rect 13820 12180 13872 12232
rect 15016 12180 15068 12232
rect 15844 12180 15896 12232
rect 5908 12112 5960 12164
rect 7104 12112 7156 12164
rect 7932 12112 7984 12164
rect 8208 12112 8260 12164
rect 9404 12112 9456 12164
rect 4068 12044 4120 12096
rect 6552 12044 6604 12096
rect 8300 12044 8352 12096
rect 9312 12087 9364 12096
rect 9312 12053 9321 12087
rect 9321 12053 9355 12087
rect 9355 12053 9364 12087
rect 9312 12044 9364 12053
rect 3566 11942 3618 11994
rect 3630 11942 3682 11994
rect 3694 11942 3746 11994
rect 3758 11942 3810 11994
rect 3822 11942 3874 11994
rect 8566 11942 8618 11994
rect 8630 11942 8682 11994
rect 8694 11942 8746 11994
rect 8758 11942 8810 11994
rect 8822 11942 8874 11994
rect 13820 11908 13872 11960
rect 15476 11908 15528 11960
rect 7564 11840 7616 11892
rect 9036 11840 9088 11892
rect 3056 11772 3108 11824
rect 5816 11815 5868 11824
rect 5816 11781 5825 11815
rect 5825 11781 5859 11815
rect 5859 11781 5868 11815
rect 5816 11772 5868 11781
rect 7104 11772 7156 11824
rect 13544 11772 13596 11824
rect 13820 11772 13872 11824
rect 16488 11772 16540 11824
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 8944 11704 8996 11756
rect 3240 11636 3292 11688
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 3608 11636 3660 11645
rect 4160 11679 4212 11688
rect 4160 11645 4169 11679
rect 4169 11645 4203 11679
rect 4203 11645 4212 11679
rect 4160 11636 4212 11645
rect 6368 11679 6420 11688
rect 6368 11645 6377 11679
rect 6377 11645 6411 11679
rect 6411 11645 6420 11679
rect 6368 11636 6420 11645
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 1860 11543 1912 11552
rect 1860 11509 1869 11543
rect 1869 11509 1903 11543
rect 1903 11509 1912 11543
rect 1860 11500 1912 11509
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 7566 11398 7618 11450
rect 7630 11398 7682 11450
rect 7694 11398 7746 11450
rect 7758 11398 7810 11450
rect 7822 11398 7874 11450
rect 13544 11432 13596 11484
rect 15660 11432 15712 11484
rect 2136 11339 2188 11348
rect 2136 11305 2145 11339
rect 2145 11305 2179 11339
rect 2179 11305 2188 11339
rect 2136 11296 2188 11305
rect 2688 11203 2740 11212
rect 2688 11169 2697 11203
rect 2697 11169 2731 11203
rect 2731 11169 2740 11203
rect 2688 11160 2740 11169
rect 4620 11160 4672 11212
rect 1860 11092 1912 11144
rect 5816 11092 5868 11144
rect 8484 11092 8536 11144
rect 3240 11067 3292 11076
rect 3240 11033 3249 11067
rect 3249 11033 3283 11067
rect 3283 11033 3292 11067
rect 3240 11024 3292 11033
rect 5540 11067 5592 11076
rect 5540 11033 5549 11067
rect 5549 11033 5583 11067
rect 5583 11033 5592 11067
rect 5540 11024 5592 11033
rect 7196 11067 7248 11076
rect 7196 11033 7205 11067
rect 7205 11033 7239 11067
rect 7239 11033 7248 11067
rect 7196 11024 7248 11033
rect 7472 11024 7524 11076
rect 4068 10956 4120 11008
rect 5172 10956 5224 11008
rect 5632 10956 5684 11008
rect 8208 11024 8260 11076
rect 14832 11024 14884 11076
rect 18144 11024 18196 11076
rect 14096 10956 14148 11008
rect 3566 10854 3618 10906
rect 3630 10854 3682 10906
rect 3694 10854 3746 10906
rect 3758 10854 3810 10906
rect 3822 10854 3874 10906
rect 8566 10854 8618 10906
rect 8630 10854 8682 10906
rect 8694 10854 8746 10906
rect 8758 10854 8810 10906
rect 8822 10854 8874 10906
rect 4804 10795 4856 10804
rect 4804 10761 4813 10795
rect 4813 10761 4847 10795
rect 4847 10761 4856 10795
rect 4804 10752 4856 10761
rect 3884 10684 3936 10736
rect 5724 10684 5776 10736
rect 7196 10684 7248 10736
rect 1676 10616 1728 10668
rect 2136 10616 2188 10668
rect 4344 10659 4396 10668
rect 4344 10625 4353 10659
rect 4353 10625 4387 10659
rect 4387 10625 4396 10659
rect 4344 10616 4396 10625
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 6184 10616 6236 10668
rect 8300 10659 8352 10668
rect 8300 10625 8309 10659
rect 8309 10625 8343 10659
rect 8343 10625 8352 10659
rect 8300 10616 8352 10625
rect 8392 10616 8444 10668
rect 2504 10591 2556 10600
rect 2504 10557 2513 10591
rect 2513 10557 2547 10591
rect 2547 10557 2556 10591
rect 2504 10548 2556 10557
rect 6736 10480 6788 10532
rect 13820 10480 13872 10532
rect 16948 10480 17000 10532
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 6276 10412 6328 10464
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 7566 10310 7618 10362
rect 7630 10310 7682 10362
rect 7694 10310 7746 10362
rect 7758 10310 7810 10362
rect 7822 10310 7874 10362
rect 13820 10276 13872 10328
rect 18420 10276 18472 10328
rect 2136 10251 2188 10260
rect 2136 10217 2145 10251
rect 2145 10217 2179 10251
rect 2179 10217 2188 10251
rect 2136 10208 2188 10217
rect 8944 10251 8996 10260
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 13728 10140 13780 10192
rect 18420 10140 18472 10192
rect 1492 10115 1544 10124
rect 1492 10081 1501 10115
rect 1501 10081 1535 10115
rect 1535 10081 1544 10115
rect 1492 10072 1544 10081
rect 2320 10072 2372 10124
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 9680 10072 9732 10124
rect 10508 10072 10560 10124
rect 15568 10072 15620 10124
rect 3424 10004 3476 10056
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 8116 10004 8168 10056
rect 5448 9936 5500 9988
rect 7012 9936 7064 9988
rect 9312 9979 9364 9988
rect 9312 9945 9321 9979
rect 9321 9945 9355 9979
rect 9355 9945 9364 9979
rect 9312 9936 9364 9945
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 3884 9868 3936 9920
rect 4068 9868 4120 9920
rect 6644 9868 6696 9920
rect 6828 9868 6880 9920
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 8300 9868 8352 9920
rect 13912 9868 13964 9920
rect 14096 9868 14148 9920
rect 15476 9868 15528 9920
rect 3566 9766 3618 9818
rect 3630 9766 3682 9818
rect 3694 9766 3746 9818
rect 3758 9766 3810 9818
rect 3822 9766 3874 9818
rect 8566 9766 8618 9818
rect 8630 9766 8682 9818
rect 8694 9766 8746 9818
rect 8758 9766 8810 9818
rect 8822 9766 8874 9818
rect 4620 9596 4672 9648
rect 9312 9664 9364 9716
rect 7380 9639 7432 9648
rect 7380 9605 7389 9639
rect 7389 9605 7423 9639
rect 7423 9605 7432 9639
rect 7380 9596 7432 9605
rect 15292 9596 15344 9648
rect 3240 9528 3292 9580
rect 3976 9528 4028 9580
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 6460 9571 6512 9580
rect 6460 9537 6469 9571
rect 6469 9537 6503 9571
rect 6503 9537 6512 9571
rect 6460 9528 6512 9537
rect 2136 9460 2188 9512
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 2964 9460 3016 9512
rect 5816 9503 5868 9512
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 5816 9460 5868 9469
rect 13176 9460 13228 9512
rect 18052 9460 18104 9512
rect 4988 9392 5040 9444
rect 9036 9324 9088 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 7566 9222 7618 9274
rect 7630 9222 7682 9274
rect 7694 9222 7746 9274
rect 7758 9222 7810 9274
rect 7822 9222 7874 9274
rect 13820 9188 13872 9240
rect 15476 9188 15528 9240
rect 4712 9163 4764 9172
rect 4712 9129 4721 9163
rect 4721 9129 4755 9163
rect 4755 9129 4764 9163
rect 4712 9120 4764 9129
rect 1492 9052 1544 9104
rect 13820 9052 13872 9104
rect 15752 9052 15804 9104
rect 3148 8984 3200 9036
rect 7104 8984 7156 9036
rect 14280 8984 14332 9036
rect 15384 8984 15436 9036
rect 1492 8959 1544 8968
rect 1492 8925 1501 8959
rect 1501 8925 1535 8959
rect 1535 8925 1544 8959
rect 1492 8916 1544 8925
rect 4160 8916 4212 8968
rect 5448 8916 5500 8968
rect 7288 8916 7340 8968
rect 9036 8959 9088 8968
rect 9036 8925 9045 8959
rect 9045 8925 9079 8959
rect 9079 8925 9088 8959
rect 9036 8916 9088 8925
rect 13084 8916 13136 8968
rect 17684 8916 17736 8968
rect 2320 8848 2372 8900
rect 15384 8848 15436 8900
rect 15936 8848 15988 8900
rect 1768 8780 1820 8832
rect 4896 8780 4948 8832
rect 9128 8823 9180 8832
rect 9128 8789 9137 8823
rect 9137 8789 9171 8823
rect 9171 8789 9180 8823
rect 9128 8780 9180 8789
rect 3566 8678 3618 8730
rect 3630 8678 3682 8730
rect 3694 8678 3746 8730
rect 3758 8678 3810 8730
rect 3822 8678 3874 8730
rect 8566 8678 8618 8730
rect 8630 8678 8682 8730
rect 8694 8678 8746 8730
rect 8758 8678 8810 8730
rect 8822 8678 8874 8730
rect 4988 8576 5040 8628
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 5632 8576 5684 8585
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 3516 8508 3568 8560
rect 9128 8551 9180 8560
rect 9128 8517 9137 8551
rect 9137 8517 9171 8551
rect 9171 8517 9180 8551
rect 9128 8508 9180 8517
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 4436 8440 4488 8492
rect 6000 8440 6052 8492
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 11244 8440 11296 8492
rect 15200 8440 15252 8492
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 8208 8415 8260 8424
rect 2780 8372 2832 8381
rect 8208 8381 8217 8415
rect 8217 8381 8251 8415
rect 8251 8381 8260 8415
rect 8208 8372 8260 8381
rect 9588 8372 9640 8424
rect 6460 8304 6512 8356
rect 7104 8304 7156 8356
rect 13544 8304 13596 8356
rect 18512 8304 18564 8356
rect 13268 8236 13320 8288
rect 16028 8236 16080 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 7566 8134 7618 8186
rect 7630 8134 7682 8186
rect 7694 8134 7746 8186
rect 7758 8134 7810 8186
rect 7822 8134 7874 8186
rect 3884 7939 3936 7948
rect 3884 7905 3893 7939
rect 3893 7905 3927 7939
rect 3927 7905 3936 7939
rect 3884 7896 3936 7905
rect 1400 7828 1452 7880
rect 7380 7828 7432 7880
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 8484 7828 8536 7880
rect 9496 7828 9548 7880
rect 3240 7803 3292 7812
rect 3240 7769 3249 7803
rect 3249 7769 3283 7803
rect 3283 7769 3292 7803
rect 3240 7760 3292 7769
rect 5264 7803 5316 7812
rect 5264 7769 5273 7803
rect 5273 7769 5307 7803
rect 5307 7769 5316 7803
rect 5264 7760 5316 7769
rect 9220 7760 9272 7812
rect 4436 7735 4488 7744
rect 4436 7701 4445 7735
rect 4445 7701 4479 7735
rect 4479 7701 4488 7735
rect 4436 7692 4488 7701
rect 7012 7692 7064 7744
rect 9864 7692 9916 7744
rect 3566 7590 3618 7642
rect 3630 7590 3682 7642
rect 3694 7590 3746 7642
rect 3758 7590 3810 7642
rect 3822 7590 3874 7642
rect 8566 7590 8618 7642
rect 8630 7590 8682 7642
rect 8694 7590 8746 7642
rect 8758 7590 8810 7642
rect 8822 7590 8874 7642
rect 11336 7624 11388 7676
rect 15844 7624 15896 7676
rect 5632 7488 5684 7540
rect 8024 7488 8076 7540
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 1492 7420 1544 7472
rect 3424 7420 3476 7472
rect 4068 7420 4120 7472
rect 4252 7420 4304 7472
rect 4804 7420 4856 7472
rect 7104 7420 7156 7472
rect 13820 7420 13872 7472
rect 18052 7420 18104 7472
rect 8024 7352 8076 7404
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 3424 7284 3476 7336
rect 6368 7327 6420 7336
rect 6368 7293 6377 7327
rect 6377 7293 6411 7327
rect 6411 7293 6420 7327
rect 6368 7284 6420 7293
rect 6920 7284 6972 7336
rect 8944 7148 8996 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 7566 7046 7618 7098
rect 7630 7046 7682 7098
rect 7694 7046 7746 7098
rect 7758 7046 7810 7098
rect 7822 7046 7874 7098
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 2320 6808 2372 6860
rect 204 6740 256 6792
rect 1400 6740 1452 6792
rect 4252 6876 4304 6928
rect 4804 6808 4856 6860
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 6092 6783 6144 6792
rect 5632 6740 5684 6749
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 7472 6740 7524 6792
rect 9036 6740 9088 6792
rect 9220 6740 9272 6792
rect 13820 6740 13872 6792
rect 15660 6740 15712 6792
rect 4804 6672 4856 6724
rect 7104 6672 7156 6724
rect 3148 6604 3200 6656
rect 5540 6604 5592 6656
rect 8484 6604 8536 6656
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 3566 6502 3618 6554
rect 3630 6502 3682 6554
rect 3694 6502 3746 6554
rect 3758 6502 3810 6554
rect 3822 6502 3874 6554
rect 8566 6502 8618 6554
rect 8630 6502 8682 6554
rect 8694 6502 8746 6554
rect 8758 6502 8810 6554
rect 8822 6502 8874 6554
rect 2688 6400 2740 6452
rect 3056 6400 3108 6452
rect 3424 6400 3476 6452
rect 4804 6332 4856 6384
rect 5632 6400 5684 6452
rect 7380 6332 7432 6384
rect 6276 6264 6328 6316
rect 7012 6264 7064 6316
rect 9496 6264 9548 6316
rect 3148 6196 3200 6248
rect 5448 6196 5500 6248
rect 6828 6196 6880 6248
rect 17914 6128 17966 6180
rect 18604 6128 18656 6180
rect 8116 6060 8168 6112
rect 9128 6060 9180 6112
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 7566 5958 7618 6010
rect 7630 5958 7682 6010
rect 7694 5958 7746 6010
rect 7758 5958 7810 6010
rect 7822 5958 7874 6010
rect 2228 5856 2280 5908
rect 2964 5856 3016 5908
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 6920 5856 6972 5908
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 388 5788 440 5840
rect 2688 5788 2740 5840
rect 3424 5720 3476 5772
rect 4804 5720 4856 5772
rect 6552 5788 6604 5840
rect 9220 5788 9272 5840
rect 13820 5788 13872 5840
rect 15568 5788 15620 5840
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 3516 5652 3568 5704
rect 8116 5720 8168 5772
rect 9036 5720 9088 5772
rect 19064 5720 19116 5772
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 1676 5584 1728 5636
rect 3148 5584 3200 5636
rect 7932 5584 7984 5636
rect 8852 5584 8904 5636
rect 10048 5584 10100 5636
rect 13820 5584 13872 5636
rect 19064 5584 19116 5636
rect 2688 5516 2740 5568
rect 9036 5559 9088 5568
rect 9036 5525 9045 5559
rect 9045 5525 9079 5559
rect 9079 5525 9088 5559
rect 9036 5516 9088 5525
rect 13728 5516 13780 5568
rect 14188 5516 14240 5568
rect 3566 5414 3618 5466
rect 3630 5414 3682 5466
rect 3694 5414 3746 5466
rect 3758 5414 3810 5466
rect 3822 5414 3874 5466
rect 8566 5414 8618 5466
rect 8630 5414 8682 5466
rect 8694 5414 8746 5466
rect 8758 5414 8810 5466
rect 8822 5414 8874 5466
rect 112 5312 164 5364
rect 2504 5312 2556 5364
rect 4068 5355 4120 5364
rect 4068 5321 4077 5355
rect 4077 5321 4111 5355
rect 4111 5321 4120 5355
rect 4068 5312 4120 5321
rect 6460 5312 6512 5364
rect 6920 5312 6972 5364
rect 8208 5312 8260 5364
rect 9956 5312 10008 5364
rect 664 5244 716 5296
rect 2320 5244 2372 5296
rect 4896 5244 4948 5296
rect 6552 5287 6604 5296
rect 6552 5253 6561 5287
rect 6561 5253 6595 5287
rect 6595 5253 6604 5287
rect 6552 5244 6604 5253
rect 6736 5244 6788 5296
rect 8576 5244 8628 5296
rect 9220 5287 9272 5296
rect 9220 5253 9229 5287
rect 9229 5253 9263 5287
rect 9263 5253 9272 5287
rect 9220 5244 9272 5253
rect 13636 5244 13688 5296
rect 17132 5244 17184 5296
rect 5264 5176 5316 5228
rect 4252 5108 4304 5160
rect 6828 5108 6880 5160
rect 8208 5176 8260 5228
rect 9772 5176 9824 5228
rect 6644 4972 6696 5024
rect 7566 4870 7618 4922
rect 7630 4870 7682 4922
rect 7694 4870 7746 4922
rect 7758 4870 7810 4922
rect 7822 4870 7874 4922
rect 3976 4768 4028 4820
rect 4712 4811 4764 4820
rect 4712 4777 4721 4811
rect 4721 4777 4755 4811
rect 4755 4777 4764 4811
rect 4712 4768 4764 4777
rect 5356 4768 5408 4820
rect 6092 4768 6144 4820
rect 7380 4811 7432 4820
rect 7380 4777 7389 4811
rect 7389 4777 7423 4811
rect 7423 4777 7432 4811
rect 7380 4768 7432 4777
rect 8300 4768 8352 4820
rect 9404 4768 9456 4820
rect 12348 4768 12400 4820
rect 17408 4768 17460 4820
rect 480 4700 532 4752
rect 5540 4700 5592 4752
rect 2044 4632 2096 4684
rect 2596 4632 2648 4684
rect 1216 4564 1268 4616
rect 2872 4564 2924 4616
rect 3516 4607 3568 4616
rect 3516 4573 3525 4607
rect 3525 4573 3559 4607
rect 3559 4573 3568 4607
rect 3516 4564 3568 4573
rect 4528 4607 4580 4616
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 4896 4564 4948 4616
rect 5448 4564 5500 4616
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 8116 4632 8168 4684
rect 7380 4564 7432 4616
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 9680 4564 9732 4616
rect 848 4496 900 4548
rect 2964 4496 3016 4548
rect 6736 4428 6788 4480
rect 3566 4326 3618 4378
rect 3630 4326 3682 4378
rect 3694 4326 3746 4378
rect 3758 4326 3810 4378
rect 3822 4326 3874 4378
rect 8566 4326 8618 4378
rect 8630 4326 8682 4378
rect 8694 4326 8746 4378
rect 8758 4326 8810 4378
rect 8822 4326 8874 4378
rect 3516 4224 3568 4276
rect 5724 4224 5776 4276
rect 7104 4224 7156 4276
rect 7380 4224 7432 4276
rect 10876 4224 10928 4276
rect 18236 4224 18288 4276
rect 3424 4156 3476 4208
rect 2688 4088 2740 4140
rect 6460 4156 6512 4208
rect 4896 4088 4948 4140
rect 5540 4088 5592 4140
rect 6092 4131 6144 4140
rect 6092 4097 6101 4131
rect 6101 4097 6135 4131
rect 6135 4097 6144 4131
rect 6092 4088 6144 4097
rect 6276 4131 6328 4140
rect 6276 4097 6285 4131
rect 6285 4097 6319 4131
rect 6319 4097 6328 4131
rect 6276 4088 6328 4097
rect 6552 4088 6604 4140
rect 4068 4063 4120 4072
rect 4068 4029 4077 4063
rect 4077 4029 4111 4063
rect 4111 4029 4120 4063
rect 4068 4020 4120 4029
rect 5816 4020 5868 4072
rect 8484 4088 8536 4140
rect 4988 3952 5040 4004
rect 6276 3952 6328 4004
rect 10784 3952 10836 4004
rect 4068 3884 4120 3936
rect 4712 3884 4764 3936
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 13820 3884 13872 3936
rect 16856 3884 16908 3936
rect 7566 3782 7618 3834
rect 7630 3782 7682 3834
rect 7694 3782 7746 3834
rect 7758 3782 7810 3834
rect 7822 3782 7874 3834
rect 3056 3680 3108 3732
rect 4620 3680 4672 3732
rect 5080 3680 5132 3732
rect 6000 3723 6052 3732
rect 6000 3689 6009 3723
rect 6009 3689 6043 3723
rect 6043 3689 6052 3723
rect 6000 3680 6052 3689
rect 2964 3476 3016 3528
rect 4712 3544 4764 3596
rect 6184 3544 6236 3596
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 6920 3476 6972 3528
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 8300 3544 8352 3596
rect 9956 3544 10008 3596
rect 7012 3476 7064 3485
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 8944 3476 8996 3528
rect 7932 3408 7984 3460
rect 11796 3408 11848 3460
rect 12256 3408 12308 3460
rect 12900 3408 12952 3460
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 8116 3340 8168 3392
rect 9220 3383 9272 3392
rect 9220 3349 9229 3383
rect 9229 3349 9263 3383
rect 9263 3349 9272 3383
rect 9220 3340 9272 3349
rect 3566 3238 3618 3290
rect 3630 3238 3682 3290
rect 3694 3238 3746 3290
rect 3758 3238 3810 3290
rect 3822 3238 3874 3290
rect 8566 3238 8618 3290
rect 8630 3238 8682 3290
rect 8694 3238 8746 3290
rect 8758 3238 8810 3290
rect 8822 3238 8874 3290
rect 5264 3136 5316 3188
rect 6276 3136 6328 3188
rect 7472 3136 7524 3188
rect 8024 3136 8076 3188
rect 3976 3111 4028 3120
rect 3976 3077 3985 3111
rect 3985 3077 4019 3111
rect 4019 3077 4028 3111
rect 3976 3068 4028 3077
rect 6644 3068 6696 3120
rect 2872 3000 2924 3052
rect 3700 3000 3752 3052
rect 4712 3043 4764 3052
rect 4712 3009 4721 3043
rect 4721 3009 4755 3043
rect 4755 3009 4764 3043
rect 4712 3000 4764 3009
rect 5172 3000 5224 3052
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 6368 3000 6420 3052
rect 6552 2932 6604 2984
rect 9864 3136 9916 3188
rect 10048 3068 10100 3120
rect 7840 2864 7892 2916
rect 9036 3000 9088 3052
rect 8576 2932 8628 2984
rect 9220 2907 9272 2916
rect 9220 2873 9229 2907
rect 9229 2873 9263 2907
rect 9263 2873 9272 2907
rect 9220 2864 9272 2873
rect 5540 2796 5592 2848
rect 8208 2796 8260 2848
rect 7566 2694 7618 2746
rect 7630 2694 7682 2746
rect 7694 2694 7746 2746
rect 7758 2694 7810 2746
rect 7822 2694 7874 2746
rect 17592 2728 17644 2780
rect 17960 2728 18012 2780
rect 3976 2592 4028 2644
rect 8576 2635 8628 2644
rect 8576 2601 8585 2635
rect 8585 2601 8619 2635
rect 8619 2601 8628 2635
rect 8576 2592 8628 2601
rect 9404 2592 9456 2644
rect 5632 2524 5684 2576
rect 5540 2456 5592 2508
rect 2780 2388 2832 2440
rect 3700 2431 3752 2440
rect 3700 2397 3709 2431
rect 3709 2397 3743 2431
rect 3743 2397 3752 2431
rect 3700 2388 3752 2397
rect 5908 2431 5960 2440
rect 5908 2397 5917 2431
rect 5917 2397 5951 2431
rect 5951 2397 5960 2431
rect 5908 2388 5960 2397
rect 6276 2388 6328 2440
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 8208 2388 8260 2440
rect 9128 2388 9180 2440
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 8300 2320 8352 2372
rect 4712 2295 4764 2304
rect 4712 2261 4721 2295
rect 4721 2261 4755 2295
rect 4755 2261 4764 2295
rect 4712 2252 4764 2261
rect 6000 2295 6052 2304
rect 6000 2261 6009 2295
rect 6009 2261 6043 2295
rect 6043 2261 6052 2295
rect 6000 2252 6052 2261
rect 6736 2295 6788 2304
rect 6736 2261 6745 2295
rect 6745 2261 6779 2295
rect 6779 2261 6788 2295
rect 6736 2252 6788 2261
rect 6828 2252 6880 2304
rect 3566 2150 3618 2202
rect 3630 2150 3682 2202
rect 3694 2150 3746 2202
rect 3758 2150 3810 2202
rect 3822 2150 3874 2202
rect 8566 2150 8618 2202
rect 8630 2150 8682 2202
rect 8694 2150 8746 2202
rect 8758 2150 8810 2202
rect 8822 2150 8874 2202
rect 4068 2048 4120 2100
rect 4344 2091 4396 2100
rect 4344 2057 4353 2091
rect 4353 2057 4387 2091
rect 4387 2057 4396 2091
rect 4344 2048 4396 2057
rect 5356 2048 5408 2100
rect 5632 2091 5684 2100
rect 5632 2057 5641 2091
rect 5641 2057 5675 2091
rect 5675 2057 5684 2091
rect 5632 2048 5684 2057
rect 6644 2048 6696 2100
rect 8944 2048 8996 2100
rect 9220 2091 9272 2100
rect 9220 2057 9229 2091
rect 9229 2057 9263 2091
rect 9263 2057 9272 2091
rect 9220 2048 9272 2057
rect 3424 1912 3476 1964
rect 4160 1955 4212 1964
rect 4160 1921 4169 1955
rect 4169 1921 4203 1955
rect 4203 1921 4212 1955
rect 4160 1912 4212 1921
rect 4804 1955 4856 1964
rect 4804 1921 4813 1955
rect 4813 1921 4847 1955
rect 4847 1921 4856 1955
rect 4804 1912 4856 1921
rect 5448 1955 5500 1964
rect 5448 1921 5457 1955
rect 5457 1921 5491 1955
rect 5491 1921 5500 1955
rect 5448 1912 5500 1921
rect 6092 1955 6144 1964
rect 6092 1921 6101 1955
rect 6101 1921 6135 1955
rect 6135 1921 6144 1955
rect 6092 1912 6144 1921
rect 6276 1955 6328 1964
rect 6276 1921 6285 1955
rect 6285 1921 6319 1955
rect 6319 1921 6328 1955
rect 6276 1912 6328 1921
rect 6828 1912 6880 1964
rect 8116 1980 8168 2032
rect 7012 1912 7064 1964
rect 9036 1912 9088 1964
rect 9312 1955 9364 1964
rect 9312 1921 9321 1955
rect 9321 1921 9355 1955
rect 9355 1921 9364 1955
rect 9312 1912 9364 1921
rect 7472 1819 7524 1828
rect 7472 1785 7481 1819
rect 7481 1785 7515 1819
rect 7515 1785 7524 1819
rect 7472 1776 7524 1785
rect 6184 1751 6236 1760
rect 6184 1717 6193 1751
rect 6193 1717 6227 1751
rect 6227 1717 6236 1751
rect 6184 1708 6236 1717
rect 7566 1606 7618 1658
rect 7630 1606 7682 1658
rect 7694 1606 7746 1658
rect 7758 1606 7810 1658
rect 7822 1606 7874 1658
rect 756 1504 808 1556
rect 4804 1504 4856 1556
rect 6552 1504 6604 1556
rect 4528 1368 4580 1420
rect 3608 1343 3660 1352
rect 3608 1309 3617 1343
rect 3617 1309 3651 1343
rect 3651 1309 3660 1343
rect 3608 1300 3660 1309
rect 4160 1343 4212 1352
rect 3240 1232 3292 1284
rect 4160 1309 4169 1343
rect 4169 1309 4203 1343
rect 4203 1309 4212 1343
rect 4160 1300 4212 1309
rect 5080 1300 5132 1352
rect 6276 1300 6328 1352
rect 6736 1343 6788 1352
rect 6736 1309 6745 1343
rect 6745 1309 6779 1343
rect 6779 1309 6788 1343
rect 6736 1300 6788 1309
rect 7380 1343 7432 1352
rect 7380 1309 7389 1343
rect 7389 1309 7423 1343
rect 7423 1309 7432 1343
rect 7380 1300 7432 1309
rect 4068 1232 4120 1284
rect 8208 1232 8260 1284
rect 4344 1207 4396 1216
rect 4344 1173 4353 1207
rect 4353 1173 4387 1207
rect 4387 1173 4396 1207
rect 4344 1164 4396 1173
rect 4896 1207 4948 1216
rect 4896 1173 4905 1207
rect 4905 1173 4939 1207
rect 4939 1173 4948 1207
rect 4896 1164 4948 1173
rect 6000 1207 6052 1216
rect 6000 1173 6009 1207
rect 6009 1173 6043 1207
rect 6043 1173 6052 1207
rect 6000 1164 6052 1173
rect 3566 1062 3618 1114
rect 3630 1062 3682 1114
rect 3694 1062 3746 1114
rect 3758 1062 3810 1114
rect 3822 1062 3874 1114
rect 8566 1062 8618 1114
rect 8630 1062 8682 1114
rect 8694 1062 8746 1114
rect 8758 1062 8810 1114
rect 8822 1062 8874 1114
<< metal2 >>
rect 938 16200 994 17000
rect 1398 16200 1454 17000
rect 1858 16200 1914 17000
rect 2318 16200 2374 17000
rect 2410 16960 2466 16969
rect 2410 16895 2466 16904
rect 386 15328 442 15337
rect 386 15263 442 15272
rect 296 14816 348 14822
rect 296 14758 348 14764
rect 202 14512 258 14521
rect 202 14447 258 14456
rect 112 13388 164 13394
rect 112 13330 164 13336
rect 124 5370 152 13330
rect 216 6798 244 14447
rect 204 6792 256 6798
rect 204 6734 256 6740
rect 112 5364 164 5370
rect 112 5306 164 5312
rect 308 1601 336 14758
rect 400 5846 428 15263
rect 952 15094 980 16200
rect 1124 15428 1176 15434
rect 1124 15370 1176 15376
rect 940 15088 992 15094
rect 940 15030 992 15036
rect 478 14920 534 14929
rect 478 14855 534 14864
rect 388 5840 440 5846
rect 388 5782 440 5788
rect 492 4758 520 14855
rect 848 12640 900 12646
rect 848 12582 900 12588
rect 664 12436 716 12442
rect 664 12378 716 12384
rect 570 12200 626 12209
rect 570 12135 626 12144
rect 480 4752 532 4758
rect 480 4694 532 4700
rect 294 1592 350 1601
rect 294 1527 350 1536
rect 584 1193 612 12135
rect 676 5302 704 12378
rect 754 9752 810 9761
rect 754 9687 810 9696
rect 664 5296 716 5302
rect 664 5238 716 5244
rect 768 1562 796 9687
rect 860 4554 888 12582
rect 938 11112 994 11121
rect 938 11047 994 11056
rect 848 4548 900 4554
rect 848 4490 900 4496
rect 756 1556 808 1562
rect 756 1498 808 1504
rect 952 1465 980 11047
rect 1136 9081 1164 15370
rect 1308 15360 1360 15366
rect 1308 15302 1360 15308
rect 1214 13832 1270 13841
rect 1214 13767 1270 13776
rect 1228 12442 1256 13767
rect 1216 12436 1268 12442
rect 1216 12378 1268 12384
rect 1320 12322 1348 15302
rect 1412 14958 1440 16200
rect 1768 15496 1820 15502
rect 1766 15464 1768 15473
rect 1820 15464 1822 15473
rect 1766 15399 1822 15408
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1688 15026 1716 15098
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1596 14906 1624 14962
rect 1872 14906 1900 16200
rect 2332 15178 2360 16200
rect 2424 15706 2452 16895
rect 2778 16200 2834 17000
rect 3146 16824 3202 16833
rect 3146 16759 3202 16768
rect 2792 15994 2820 16200
rect 2792 15966 3004 15994
rect 2566 15804 2874 15813
rect 2566 15802 2572 15804
rect 2628 15802 2652 15804
rect 2708 15802 2732 15804
rect 2788 15802 2812 15804
rect 2868 15802 2874 15804
rect 2628 15750 2630 15802
rect 2810 15750 2812 15802
rect 2566 15748 2572 15750
rect 2628 15748 2652 15750
rect 2708 15748 2732 15750
rect 2788 15748 2812 15750
rect 2868 15748 2874 15750
rect 2566 15739 2874 15748
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2780 15360 2832 15366
rect 2778 15328 2780 15337
rect 2832 15328 2834 15337
rect 2778 15263 2834 15272
rect 1412 13394 1440 14894
rect 1596 14878 1900 14906
rect 2240 15150 2360 15178
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 13938 1532 14214
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1400 13388 1452 13394
rect 1400 13330 1452 13336
rect 1400 13252 1452 13258
rect 1400 13194 1452 13200
rect 1228 12294 1348 12322
rect 1122 9072 1178 9081
rect 1122 9007 1178 9016
rect 1122 8392 1178 8401
rect 1122 8327 1178 8336
rect 1030 7848 1086 7857
rect 1030 7783 1086 7792
rect 938 1456 994 1465
rect 938 1391 994 1400
rect 570 1184 626 1193
rect 570 1119 626 1128
rect 1044 921 1072 7783
rect 1136 1329 1164 8327
rect 1228 4622 1256 12294
rect 1306 12064 1362 12073
rect 1306 11999 1362 12008
rect 1320 4729 1348 11999
rect 1412 11665 1440 13194
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 12481 1624 13126
rect 1582 12472 1638 12481
rect 1582 12407 1638 12416
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1398 11656 1454 11665
rect 1398 11591 1454 11600
rect 1412 7886 1440 11591
rect 1504 10130 1532 12038
rect 1688 10674 1716 14878
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1780 12850 1808 13670
rect 2240 13297 2268 15150
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2226 13288 2282 13297
rect 2226 13223 2282 13232
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1504 9110 1532 10066
rect 1492 9104 1544 9110
rect 1492 9046 1544 9052
rect 1492 8968 1544 8974
rect 1780 8922 1808 12786
rect 2134 11792 2190 11801
rect 2134 11727 2190 11736
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11150 1900 11494
rect 2148 11354 2176 11727
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 1492 8910 1544 8916
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1504 7478 1532 8910
rect 1688 8894 1808 8922
rect 1492 7472 1544 7478
rect 1492 7414 1544 7420
rect 1504 6866 1532 7414
rect 1582 6896 1638 6905
rect 1492 6860 1544 6866
rect 1582 6831 1638 6840
rect 1492 6802 1544 6808
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 5273 1440 6734
rect 1596 5710 1624 6831
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1688 5642 1716 8894
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8498 1808 8774
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1780 6866 1808 8434
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 1398 5264 1454 5273
rect 1398 5199 1454 5208
rect 1306 4720 1362 4729
rect 2056 4690 2084 10406
rect 2148 10266 2176 10610
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2332 10130 2360 14962
rect 2778 14920 2834 14929
rect 2778 14855 2780 14864
rect 2832 14855 2834 14864
rect 2780 14826 2832 14832
rect 2566 14716 2874 14725
rect 2566 14714 2572 14716
rect 2628 14714 2652 14716
rect 2708 14714 2732 14716
rect 2788 14714 2812 14716
rect 2868 14714 2874 14716
rect 2628 14662 2630 14714
rect 2810 14662 2812 14714
rect 2566 14660 2572 14662
rect 2628 14660 2652 14662
rect 2708 14660 2732 14662
rect 2788 14660 2812 14662
rect 2868 14660 2874 14662
rect 2566 14651 2874 14660
rect 2504 14340 2556 14346
rect 2504 14282 2556 14288
rect 2516 13977 2544 14282
rect 2976 14090 3004 15966
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2608 14062 3004 14090
rect 2502 13968 2558 13977
rect 2412 13932 2464 13938
rect 2502 13903 2558 13912
rect 2412 13874 2464 13880
rect 2424 12306 2452 13874
rect 2608 13818 2636 14062
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2792 13841 2820 13874
rect 2516 13790 2636 13818
rect 2778 13832 2834 13841
rect 2516 13734 2544 13790
rect 2778 13767 2834 13776
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2566 13628 2874 13637
rect 2566 13626 2572 13628
rect 2628 13626 2652 13628
rect 2708 13626 2732 13628
rect 2788 13626 2812 13628
rect 2868 13626 2874 13628
rect 2628 13574 2630 13626
rect 2810 13574 2812 13626
rect 2566 13572 2572 13574
rect 2628 13572 2652 13574
rect 2708 13572 2732 13574
rect 2788 13572 2812 13574
rect 2868 13572 2874 13574
rect 2566 13563 2874 13572
rect 2976 12850 3004 13738
rect 3068 13734 3096 15438
rect 3160 15434 3188 16759
rect 3238 16200 3294 17000
rect 3436 16238 3648 16266
rect 3252 16130 3280 16200
rect 3252 16102 3372 16130
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3146 13968 3202 13977
rect 3146 13903 3202 13912
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 3160 13546 3188 13903
rect 3068 13518 3188 13546
rect 3068 13326 3096 13518
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2596 12776 2648 12782
rect 2594 12744 2596 12753
rect 2648 12744 2650 12753
rect 2594 12679 2650 12688
rect 2566 12540 2874 12549
rect 2566 12538 2572 12540
rect 2628 12538 2652 12540
rect 2708 12538 2732 12540
rect 2788 12538 2812 12540
rect 2868 12538 2874 12540
rect 2628 12486 2630 12538
rect 2810 12486 2812 12538
rect 2566 12484 2572 12486
rect 2628 12484 2652 12486
rect 2708 12484 2732 12486
rect 2788 12484 2812 12486
rect 2868 12484 2874 12486
rect 2566 12475 2874 12484
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 3068 12170 3096 13262
rect 3252 12238 3280 14350
rect 3344 13002 3372 16102
rect 3436 13433 3464 16238
rect 3620 16130 3648 16238
rect 3698 16200 3754 17000
rect 4158 16200 4214 17000
rect 4618 16200 4674 17000
rect 4710 16688 4766 16697
rect 4710 16623 4766 16632
rect 3712 16130 3740 16200
rect 3620 16102 3740 16130
rect 4066 16144 4122 16153
rect 4066 16079 4122 16088
rect 4080 15502 4108 16079
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3566 15260 3874 15269
rect 3566 15258 3572 15260
rect 3628 15258 3652 15260
rect 3708 15258 3732 15260
rect 3788 15258 3812 15260
rect 3868 15258 3874 15260
rect 3628 15206 3630 15258
rect 3810 15206 3812 15258
rect 3566 15204 3572 15206
rect 3628 15204 3652 15206
rect 3708 15204 3732 15206
rect 3788 15204 3812 15206
rect 3868 15204 3874 15206
rect 3566 15195 3874 15204
rect 4066 15056 4122 15065
rect 3516 15020 3568 15026
rect 4172 15042 4200 16200
rect 4172 15014 4384 15042
rect 4066 14991 4068 15000
rect 3516 14962 3568 14968
rect 4120 14991 4122 15000
rect 4068 14962 4120 14968
rect 3528 14346 3556 14962
rect 4080 14906 4108 14962
rect 3988 14878 4108 14906
rect 4160 14884 4212 14890
rect 3988 14550 4016 14878
rect 4160 14826 4212 14832
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 3976 14408 4028 14414
rect 3974 14376 3976 14385
rect 4028 14376 4030 14385
rect 3516 14340 3568 14346
rect 3974 14311 4030 14320
rect 3516 14282 3568 14288
rect 3976 14272 4028 14278
rect 4080 14249 4108 14758
rect 3976 14214 4028 14220
rect 4066 14240 4122 14249
rect 3566 14172 3874 14181
rect 3566 14170 3572 14172
rect 3628 14170 3652 14172
rect 3708 14170 3732 14172
rect 3788 14170 3812 14172
rect 3868 14170 3874 14172
rect 3628 14118 3630 14170
rect 3810 14118 3812 14170
rect 3566 14116 3572 14118
rect 3628 14116 3652 14118
rect 3708 14116 3732 14118
rect 3788 14116 3812 14118
rect 3868 14116 3874 14118
rect 3566 14107 3874 14116
rect 3422 13424 3478 13433
rect 3422 13359 3478 13368
rect 3566 13084 3874 13093
rect 3566 13082 3572 13084
rect 3628 13082 3652 13084
rect 3708 13082 3732 13084
rect 3788 13082 3812 13084
rect 3868 13082 3874 13084
rect 3628 13030 3630 13082
rect 3810 13030 3812 13082
rect 3566 13028 3572 13030
rect 3628 13028 3652 13030
rect 3708 13028 3732 13030
rect 3788 13028 3812 13030
rect 3868 13028 3874 13030
rect 3566 13019 3874 13028
rect 3344 12974 3464 13002
rect 3436 12434 3464 12974
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3344 12406 3464 12434
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2566 11452 2874 11461
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11387 2874 11396
rect 2686 11248 2742 11257
rect 2686 11183 2688 11192
rect 2740 11183 2742 11192
rect 2688 11154 2740 11160
rect 2504 10600 2556 10606
rect 2502 10568 2504 10577
rect 2556 10568 2558 10577
rect 2502 10503 2558 10512
rect 2566 10364 2874 10373
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10299 2874 10308
rect 2976 10169 3004 12038
rect 3068 11830 3096 12106
rect 3056 11824 3108 11830
rect 3344 11778 3372 12406
rect 3424 12232 3476 12238
rect 3528 12209 3556 12854
rect 3424 12174 3476 12180
rect 3514 12200 3570 12209
rect 3056 11766 3108 11772
rect 3160 11750 3372 11778
rect 3436 11778 3464 12174
rect 3514 12135 3570 12144
rect 3566 11996 3874 12005
rect 3566 11994 3572 11996
rect 3628 11994 3652 11996
rect 3708 11994 3732 11996
rect 3788 11994 3812 11996
rect 3868 11994 3874 11996
rect 3628 11942 3630 11994
rect 3810 11942 3812 11994
rect 3566 11940 3572 11942
rect 3628 11940 3652 11942
rect 3708 11940 3732 11942
rect 3788 11940 3812 11942
rect 3868 11940 3874 11942
rect 3566 11931 3874 11940
rect 3436 11750 3648 11778
rect 3160 11370 3188 11750
rect 3620 11694 3648 11750
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3068 11342 3188 11370
rect 2962 10160 3018 10169
rect 2320 10124 2372 10130
rect 2962 10095 3018 10104
rect 2320 10066 2372 10072
rect 2136 9512 2188 9518
rect 2688 9512 2740 9518
rect 2136 9454 2188 9460
rect 2686 9480 2688 9489
rect 2964 9512 3016 9518
rect 2740 9480 2742 9489
rect 1306 4655 1362 4664
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 1216 4616 1268 4622
rect 2148 4604 2176 9454
rect 2964 9454 3016 9460
rect 2686 9415 2742 9424
rect 2566 9276 2874 9285
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9211 2874 9220
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 2226 7440 2282 7449
rect 2226 7375 2282 7384
rect 2240 5914 2268 7375
rect 2332 6866 2360 8842
rect 2780 8424 2832 8430
rect 2778 8392 2780 8401
rect 2832 8392 2834 8401
rect 2778 8327 2834 8336
rect 2566 8188 2874 8197
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8123 2874 8132
rect 2410 7984 2466 7993
rect 2410 7919 2466 7928
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 2332 4706 2360 5238
rect 2424 4865 2452 7919
rect 2566 7100 2874 7109
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7035 2874 7044
rect 2976 6914 3004 9454
rect 3068 7993 3096 11342
rect 3252 11200 3280 11630
rect 3620 11529 3648 11630
rect 3606 11520 3662 11529
rect 3606 11455 3662 11464
rect 3160 11172 3280 11200
rect 3160 9042 3188 11172
rect 3238 11112 3294 11121
rect 3238 11047 3240 11056
rect 3292 11047 3294 11056
rect 3240 11018 3292 11024
rect 3566 10908 3874 10917
rect 3566 10906 3572 10908
rect 3628 10906 3652 10908
rect 3708 10906 3732 10908
rect 3788 10906 3812 10908
rect 3868 10906 3874 10908
rect 3628 10854 3630 10906
rect 3810 10854 3812 10906
rect 3566 10852 3572 10854
rect 3628 10852 3652 10854
rect 3708 10852 3732 10854
rect 3788 10852 3812 10854
rect 3868 10852 3874 10854
rect 3566 10843 3874 10852
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 3424 10056 3476 10062
rect 3330 10024 3386 10033
rect 3424 9998 3476 10004
rect 3330 9959 3386 9968
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3252 9761 3280 9862
rect 3238 9752 3294 9761
rect 3238 9687 3294 9696
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3054 7984 3110 7993
rect 3054 7919 3110 7928
rect 2700 6886 3004 6914
rect 3054 6896 3110 6905
rect 2700 6458 2728 6886
rect 2976 6840 3054 6848
rect 2976 6831 3110 6840
rect 2976 6820 3096 6831
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2566 6012 2874 6021
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5947 2874 5956
rect 2976 5914 3004 6820
rect 3160 6746 3188 8978
rect 3252 8945 3280 9522
rect 3238 8936 3294 8945
rect 3238 8871 3294 8880
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3252 7313 3280 7754
rect 3238 7304 3294 7313
rect 3238 7239 3294 7248
rect 3068 6718 3188 6746
rect 3068 6458 3096 6718
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 3160 6254 3188 6598
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3054 5944 3110 5953
rect 2964 5908 3016 5914
rect 3054 5879 3110 5888
rect 2964 5850 3016 5856
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2504 5704 2556 5710
rect 2502 5672 2504 5681
rect 2556 5672 2558 5681
rect 2700 5658 2728 5782
rect 2700 5630 2820 5658
rect 2502 5607 2558 5616
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2410 4856 2466 4865
rect 2410 4791 2466 4800
rect 2332 4678 2452 4706
rect 2148 4576 2360 4604
rect 1216 4558 1268 4564
rect 2332 4026 2360 4576
rect 2424 4185 2452 4678
rect 2410 4176 2466 4185
rect 2410 4111 2466 4120
rect 2410 4040 2466 4049
rect 2332 3998 2410 4026
rect 2410 3975 2466 3984
rect 2516 2689 2544 5306
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2608 3913 2636 4626
rect 2700 4146 2728 5510
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2686 4040 2742 4049
rect 2686 3975 2742 3984
rect 2594 3904 2650 3913
rect 2594 3839 2650 3848
rect 2700 3777 2728 3975
rect 2686 3768 2742 3777
rect 2686 3703 2742 3712
rect 2792 3618 2820 5630
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2700 3590 2820 3618
rect 2502 2680 2558 2689
rect 2502 2615 2558 2624
rect 2700 2553 2728 3590
rect 2884 3058 2912 4558
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2976 3534 3004 4490
rect 3068 3738 3096 5879
rect 3160 5642 3188 6190
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3146 3904 3202 3913
rect 3146 3839 3202 3848
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3160 3641 3188 3839
rect 3146 3632 3202 3641
rect 3146 3567 3202 3576
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2686 2544 2742 2553
rect 2686 2479 2742 2488
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 1858 1592 1914 1601
rect 2318 1592 2374 1601
rect 1914 1550 2318 1578
rect 1858 1527 1914 1536
rect 2318 1527 2374 1536
rect 2792 1465 2820 2382
rect 2870 1728 2926 1737
rect 2870 1663 2926 1672
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 1122 1320 1178 1329
rect 1122 1255 1178 1264
rect 2884 1193 2912 1663
rect 3252 1290 3280 7239
rect 3344 3913 3372 9959
rect 3436 7478 3464 9998
rect 3896 9926 3924 10678
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3566 9820 3874 9829
rect 3566 9818 3572 9820
rect 3628 9818 3652 9820
rect 3708 9818 3732 9820
rect 3788 9818 3812 9820
rect 3868 9818 3874 9820
rect 3628 9766 3630 9818
rect 3810 9766 3812 9818
rect 3566 9764 3572 9766
rect 3628 9764 3652 9766
rect 3708 9764 3732 9766
rect 3788 9764 3812 9766
rect 3868 9764 3874 9766
rect 3566 9755 3874 9764
rect 3988 9586 4016 14214
rect 4066 14175 4122 14184
rect 4066 14104 4122 14113
rect 4066 14039 4122 14048
rect 4080 14006 4108 14039
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4080 13161 4108 13262
rect 4066 13152 4122 13161
rect 4066 13087 4122 13096
rect 4172 12458 4200 14826
rect 4080 12430 4200 12458
rect 4080 12238 4108 12430
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4080 11121 4108 12038
rect 4160 11688 4212 11694
rect 4158 11656 4160 11665
rect 4212 11656 4214 11665
rect 4158 11591 4214 11600
rect 4066 11112 4122 11121
rect 4066 11047 4122 11056
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10130 4108 10950
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 4080 9217 4108 9862
rect 4264 9738 4292 12174
rect 4356 11937 4384 15014
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4436 14544 4488 14550
rect 4434 14512 4436 14521
rect 4488 14512 4490 14521
rect 4434 14447 4490 14456
rect 4540 13938 4568 14758
rect 4632 14498 4660 16200
rect 4724 15570 4752 16623
rect 5078 16200 5134 17000
rect 5538 16200 5594 17000
rect 5998 16200 6054 17000
rect 6182 16280 6238 16289
rect 6182 16215 6238 16224
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4632 14470 4752 14498
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4434 13016 4490 13025
rect 4434 12951 4490 12960
rect 4448 12850 4476 12951
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 4342 11928 4398 11937
rect 4342 11863 4398 11872
rect 4632 11218 4660 14470
rect 4724 14414 4752 14470
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 5092 14006 5120 16200
rect 5448 15496 5500 15502
rect 5262 15464 5318 15473
rect 5448 15438 5500 15444
rect 5552 15450 5580 16200
rect 5722 16008 5778 16017
rect 5722 15943 5778 15952
rect 5736 15706 5764 15943
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5262 15399 5318 15408
rect 5276 14482 5304 15399
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5460 15314 5488 15438
rect 5552 15422 5764 15450
rect 5368 15065 5396 15302
rect 5460 15286 5580 15314
rect 5552 15162 5580 15286
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5354 15056 5410 15065
rect 5354 14991 5410 15000
rect 5736 14958 5764 15422
rect 5724 14952 5776 14958
rect 5446 14920 5502 14929
rect 5724 14894 5776 14900
rect 5446 14855 5502 14864
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5080 14000 5132 14006
rect 4894 13968 4950 13977
rect 5080 13942 5132 13948
rect 4894 13903 4896 13912
rect 4948 13903 4950 13912
rect 4896 13874 4948 13880
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 12434 4936 12582
rect 5184 12434 5212 13262
rect 5276 12850 5304 14418
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5368 13920 5396 14282
rect 5460 14074 5488 14855
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5448 13932 5500 13938
rect 5368 13892 5448 13920
rect 5448 13874 5500 13880
rect 5460 13394 5488 13874
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 4908 12406 5028 12434
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4356 10033 4384 10610
rect 4342 10024 4398 10033
rect 4342 9959 4398 9968
rect 4172 9710 4292 9738
rect 4526 9752 4582 9761
rect 4066 9208 4122 9217
rect 4066 9143 4122 9152
rect 4172 9058 4200 9710
rect 4526 9687 4582 9696
rect 3988 9030 4200 9058
rect 3566 8732 3874 8741
rect 3566 8730 3572 8732
rect 3628 8730 3652 8732
rect 3708 8730 3732 8732
rect 3788 8730 3812 8732
rect 3868 8730 3874 8732
rect 3628 8678 3630 8730
rect 3810 8678 3812 8730
rect 3566 8676 3572 8678
rect 3628 8676 3652 8678
rect 3708 8676 3732 8678
rect 3788 8676 3812 8678
rect 3868 8676 3874 8678
rect 3566 8667 3874 8676
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3528 7857 3556 8502
rect 3882 7984 3938 7993
rect 3882 7919 3884 7928
rect 3936 7919 3938 7928
rect 3884 7890 3936 7896
rect 3514 7848 3570 7857
rect 3514 7783 3570 7792
rect 3566 7644 3874 7653
rect 3566 7642 3572 7644
rect 3628 7642 3652 7644
rect 3708 7642 3732 7644
rect 3788 7642 3812 7644
rect 3868 7642 3874 7644
rect 3628 7590 3630 7642
rect 3810 7590 3812 7642
rect 3566 7588 3572 7590
rect 3628 7588 3652 7590
rect 3708 7588 3732 7590
rect 3788 7588 3812 7590
rect 3868 7588 3874 7590
rect 3566 7579 3874 7588
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3436 7342 3464 7414
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3436 6458 3464 7278
rect 3566 6556 3874 6565
rect 3566 6554 3572 6556
rect 3628 6554 3652 6556
rect 3708 6554 3732 6556
rect 3788 6554 3812 6556
rect 3868 6554 3874 6556
rect 3628 6502 3630 6554
rect 3810 6502 3812 6554
rect 3566 6500 3572 6502
rect 3628 6500 3652 6502
rect 3708 6500 3732 6502
rect 3788 6500 3812 6502
rect 3868 6500 3874 6502
rect 3566 6491 3874 6500
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3436 5778 3464 6394
rect 3514 6352 3570 6361
rect 3514 6287 3570 6296
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3528 5710 3556 6287
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3566 5468 3874 5477
rect 3566 5466 3572 5468
rect 3628 5466 3652 5468
rect 3708 5466 3732 5468
rect 3788 5466 3812 5468
rect 3868 5466 3874 5468
rect 3628 5414 3630 5466
rect 3810 5414 3812 5466
rect 3566 5412 3572 5414
rect 3628 5412 3652 5414
rect 3708 5412 3732 5414
rect 3788 5412 3812 5414
rect 3868 5412 3874 5414
rect 3566 5403 3874 5412
rect 3988 4826 4016 9030
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4172 7698 4200 8910
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4448 7834 4476 8434
rect 4080 7670 4200 7698
rect 4356 7806 4476 7834
rect 4080 7478 4108 7670
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4066 7032 4122 7041
rect 4066 6967 4122 6976
rect 4080 5370 4108 6967
rect 4264 6934 4292 7414
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4264 5166 4292 6870
rect 4252 5160 4304 5166
rect 4158 5128 4214 5137
rect 4252 5102 4304 5108
rect 4158 5063 4214 5072
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3514 4720 3570 4729
rect 3514 4655 3570 4664
rect 3528 4622 3556 4655
rect 3516 4616 3568 4622
rect 3436 4576 3516 4604
rect 3436 4214 3464 4576
rect 3516 4558 3568 4564
rect 3566 4380 3874 4389
rect 3566 4378 3572 4380
rect 3628 4378 3652 4380
rect 3708 4378 3732 4380
rect 3788 4378 3812 4380
rect 3868 4378 3874 4380
rect 3628 4326 3630 4378
rect 3810 4326 3812 4378
rect 3566 4324 3572 4326
rect 3628 4324 3652 4326
rect 3708 4324 3732 4326
rect 3788 4324 3812 4326
rect 3868 4324 3874 4326
rect 3566 4315 3874 4324
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3528 4026 3556 4218
rect 3974 4176 4030 4185
rect 3974 4111 4030 4120
rect 3436 3998 3556 4026
rect 3330 3904 3386 3913
rect 3330 3839 3386 3848
rect 3436 1970 3464 3998
rect 3566 3292 3874 3301
rect 3566 3290 3572 3292
rect 3628 3290 3652 3292
rect 3708 3290 3732 3292
rect 3788 3290 3812 3292
rect 3868 3290 3874 3292
rect 3628 3238 3630 3290
rect 3810 3238 3812 3290
rect 3566 3236 3572 3238
rect 3628 3236 3652 3238
rect 3708 3236 3732 3238
rect 3788 3236 3812 3238
rect 3868 3236 3874 3238
rect 3566 3227 3874 3236
rect 3988 3126 4016 4111
rect 4068 4072 4120 4078
rect 4066 4040 4068 4049
rect 4120 4040 4122 4049
rect 4066 3975 4122 3984
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3712 2446 3740 2994
rect 4080 2938 4108 3878
rect 4172 3534 4200 5063
rect 4356 4128 4384 7806
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4264 4100 4384 4128
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 3988 2910 4108 2938
rect 3988 2650 4016 2910
rect 4264 2774 4292 4100
rect 4342 3904 4398 3913
rect 4342 3839 4398 3848
rect 4080 2746 4292 2774
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 3566 2204 3874 2213
rect 3566 2202 3572 2204
rect 3628 2202 3652 2204
rect 3708 2202 3732 2204
rect 3788 2202 3812 2204
rect 3868 2202 3874 2204
rect 3628 2150 3630 2202
rect 3810 2150 3812 2202
rect 3566 2148 3572 2150
rect 3628 2148 3652 2150
rect 3708 2148 3732 2150
rect 3788 2148 3812 2150
rect 3868 2148 3874 2150
rect 3566 2139 3874 2148
rect 4080 2106 4108 2746
rect 4356 2106 4384 3839
rect 4448 2774 4476 7686
rect 4540 6769 4568 9687
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4526 6760 4582 6769
rect 4526 6695 4582 6704
rect 4632 5953 4660 9590
rect 4724 9178 4752 12174
rect 4894 11520 4950 11529
rect 4894 11455 4950 11464
rect 4802 10840 4858 10849
rect 4802 10775 4804 10784
rect 4856 10775 4858 10784
rect 4804 10746 4856 10752
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4908 8838 4936 11455
rect 5000 11121 5028 12406
rect 5092 12406 5212 12434
rect 4986 11112 5042 11121
rect 4986 11047 5042 11056
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 5000 9081 5028 9386
rect 4986 9072 5042 9081
rect 4986 9007 5042 9016
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4816 6866 4844 7414
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4816 6730 4844 6802
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4816 6390 4844 6666
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4618 5944 4674 5953
rect 4618 5879 4674 5888
rect 4618 5808 4674 5817
rect 4816 5778 4844 6326
rect 4618 5743 4674 5752
rect 4804 5772 4856 5778
rect 4526 5264 4582 5273
rect 4526 5199 4582 5208
rect 4540 4622 4568 5199
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4632 3738 4660 5743
rect 4804 5714 4856 5720
rect 4802 5672 4858 5681
rect 4908 5658 4936 8774
rect 5000 8634 5028 9007
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4858 5630 4936 5658
rect 4986 5672 5042 5681
rect 4802 5607 4858 5616
rect 4986 5607 5042 5616
rect 4710 5264 4766 5273
rect 4710 5199 4766 5208
rect 4724 4826 4752 5199
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4710 4720 4766 4729
rect 4710 4655 4766 4664
rect 4724 3942 4752 4655
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4724 3058 4752 3538
rect 4816 3414 4844 5607
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 4908 4865 4936 5238
rect 4894 4856 4950 4865
rect 4894 4791 4950 4800
rect 4908 4622 4936 4791
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4908 3534 4936 4082
rect 5000 4010 5028 5607
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 5092 3738 5120 12406
rect 5460 11370 5488 13330
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 11801 5580 13262
rect 5538 11792 5594 11801
rect 5538 11727 5594 11736
rect 5460 11342 5672 11370
rect 5446 11248 5502 11257
rect 5446 11183 5502 11192
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4816 3386 5120 3414
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4448 2746 4568 2774
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4344 2100 4396 2106
rect 4344 2042 4396 2048
rect 3424 1964 3476 1970
rect 3424 1906 3476 1912
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 4172 1601 4200 1906
rect 4158 1592 4214 1601
rect 4158 1527 4214 1536
rect 4540 1426 4568 2746
rect 4712 2304 4764 2310
rect 4710 2272 4712 2281
rect 4764 2272 4766 2281
rect 4710 2207 4766 2216
rect 4804 1964 4856 1970
rect 4804 1906 4856 1912
rect 4816 1562 4844 1906
rect 4804 1556 4856 1562
rect 4804 1498 4856 1504
rect 4528 1420 4580 1426
rect 4528 1362 4580 1368
rect 5092 1358 5120 3386
rect 5184 3058 5212 10950
rect 5460 9994 5488 11183
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5368 8401 5396 9522
rect 5552 9058 5580 11018
rect 5644 11014 5672 11342
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5644 10674 5672 10950
rect 5736 10742 5764 14894
rect 6012 13920 6040 16200
rect 6196 15502 6224 16215
rect 6458 16200 6514 17000
rect 18418 16960 18474 16969
rect 18418 16895 18474 16904
rect 13634 16824 13690 16833
rect 13634 16759 13690 16768
rect 13648 16726 13676 16759
rect 13636 16720 13688 16726
rect 15292 16720 15344 16726
rect 13636 16662 13688 16668
rect 13726 16688 13782 16697
rect 13726 16623 13782 16632
rect 15106 16688 15162 16697
rect 15106 16623 15162 16632
rect 15290 16688 15292 16697
rect 15344 16688 15346 16697
rect 15290 16623 15346 16632
rect 18234 16688 18290 16697
rect 18234 16623 18290 16632
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6472 14414 6500 16200
rect 13082 16144 13138 16153
rect 13082 16079 13138 16088
rect 7566 15804 7874 15813
rect 7566 15802 7572 15804
rect 7628 15802 7652 15804
rect 7708 15802 7732 15804
rect 7788 15802 7812 15804
rect 7868 15802 7874 15804
rect 7628 15750 7630 15802
rect 7810 15750 7812 15802
rect 7566 15748 7572 15750
rect 7628 15748 7652 15750
rect 7708 15748 7732 15750
rect 7788 15748 7812 15750
rect 7868 15748 7874 15750
rect 7566 15739 7874 15748
rect 8392 15496 8444 15502
rect 8114 15464 8170 15473
rect 7840 15428 7892 15434
rect 8392 15438 8444 15444
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 11058 15464 11114 15473
rect 8114 15399 8116 15408
rect 7840 15370 7892 15376
rect 8168 15399 8170 15408
rect 8116 15370 8168 15376
rect 6550 15192 6606 15201
rect 6550 15127 6606 15136
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6012 13892 6132 13920
rect 6000 13796 6052 13802
rect 6000 13738 6052 13744
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5828 11830 5856 12718
rect 6012 12209 6040 13738
rect 6104 12345 6132 13892
rect 6564 12850 6592 15127
rect 7852 15094 7880 15370
rect 8404 15201 8432 15438
rect 8566 15260 8874 15269
rect 8566 15258 8572 15260
rect 8628 15258 8652 15260
rect 8708 15258 8732 15260
rect 8788 15258 8812 15260
rect 8868 15258 8874 15260
rect 8628 15206 8630 15258
rect 8810 15206 8812 15258
rect 8566 15204 8572 15206
rect 8628 15204 8652 15206
rect 8708 15204 8732 15206
rect 8788 15204 8812 15206
rect 8868 15204 8874 15206
rect 8390 15192 8446 15201
rect 8566 15195 8874 15204
rect 8390 15127 8446 15136
rect 7840 15088 7892 15094
rect 8208 15088 8260 15094
rect 7892 15036 7972 15042
rect 7840 15030 7972 15036
rect 8208 15030 8260 15036
rect 7852 15014 7972 15030
rect 7566 14716 7874 14725
rect 7566 14714 7572 14716
rect 7628 14714 7652 14716
rect 7708 14714 7732 14716
rect 7788 14714 7812 14716
rect 7868 14714 7874 14716
rect 7628 14662 7630 14714
rect 7810 14662 7812 14714
rect 7566 14660 7572 14662
rect 7628 14660 7652 14662
rect 7708 14660 7732 14662
rect 7788 14660 7812 14662
rect 7868 14660 7874 14662
rect 7566 14651 7874 14660
rect 6918 14376 6974 14385
rect 6918 14311 6974 14320
rect 7380 14340 7432 14346
rect 6644 13864 6696 13870
rect 6642 13832 6644 13841
rect 6696 13832 6698 13841
rect 6642 13767 6698 13776
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6656 12889 6684 13194
rect 6642 12880 6698 12889
rect 6552 12844 6604 12850
rect 6642 12815 6698 12824
rect 6552 12786 6604 12792
rect 6564 12434 6592 12786
rect 6380 12406 6592 12434
rect 6090 12336 6146 12345
rect 6090 12271 6146 12280
rect 5998 12200 6054 12209
rect 5908 12164 5960 12170
rect 5998 12135 6054 12144
rect 5908 12106 5960 12112
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5644 9761 5672 10610
rect 5630 9752 5686 9761
rect 5828 9738 5856 11086
rect 5630 9687 5686 9696
rect 5736 9710 5856 9738
rect 5460 9030 5580 9058
rect 5460 8974 5488 9030
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5644 8537 5672 8570
rect 5630 8528 5686 8537
rect 5630 8463 5686 8472
rect 5354 8392 5410 8401
rect 5354 8327 5410 8336
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5276 5234 5304 7754
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5354 7168 5410 7177
rect 5354 7103 5410 7112
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5368 4826 5396 7103
rect 5644 6882 5672 7482
rect 5460 6854 5672 6882
rect 5460 6254 5488 6854
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5446 6080 5502 6089
rect 5446 6015 5502 6024
rect 5460 5001 5488 6015
rect 5552 5914 5580 6598
rect 5644 6458 5672 6734
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5446 4992 5502 5001
rect 5446 4927 5502 4936
rect 5446 4856 5502 4865
rect 5356 4820 5408 4826
rect 5446 4791 5502 4800
rect 5356 4762 5408 4768
rect 5460 4622 5488 4791
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5262 4312 5318 4321
rect 5262 4247 5318 4256
rect 5276 3194 5304 4247
rect 5552 4146 5580 4694
rect 5736 4282 5764 9710
rect 5814 9616 5870 9625
rect 5814 9551 5870 9560
rect 5828 9518 5856 9551
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5814 9208 5870 9217
rect 5814 9143 5870 9152
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5828 4078 5856 9143
rect 5920 4321 5948 12106
rect 6104 11393 6132 12271
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6288 11665 6316 12174
rect 6380 11694 6408 12406
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6368 11688 6420 11694
rect 6274 11656 6330 11665
rect 6368 11630 6420 11636
rect 6274 11591 6330 11600
rect 6380 11529 6408 11630
rect 6366 11520 6422 11529
rect 6366 11455 6422 11464
rect 6090 11384 6146 11393
rect 6090 11319 6146 11328
rect 6458 11112 6514 11121
rect 6458 11047 6514 11056
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6012 9761 6040 9998
rect 5998 9752 6054 9761
rect 5998 9687 6054 9696
rect 5998 9344 6054 9353
rect 5998 9279 6054 9288
rect 6012 8498 6040 9279
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 5998 6216 6054 6225
rect 5998 6151 6054 6160
rect 5906 4312 5962 4321
rect 5906 4247 5962 4256
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5460 3777 5488 3878
rect 5446 3768 5502 3777
rect 6012 3738 6040 6151
rect 6104 4826 6132 6734
rect 6196 5817 6224 10610
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6288 6497 6316 10406
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6380 8634 6408 9998
rect 6472 9586 6500 11047
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6380 7041 6408 7278
rect 6366 7032 6422 7041
rect 6366 6967 6422 6976
rect 6472 6882 6500 8298
rect 6380 6854 6500 6882
rect 6274 6488 6330 6497
rect 6274 6423 6330 6432
rect 6288 6322 6316 6423
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6182 5808 6238 5817
rect 6182 5743 6238 5752
rect 6380 5556 6408 6854
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6288 5528 6408 5556
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6182 4720 6238 4729
rect 6182 4655 6238 4664
rect 6196 4622 6224 4655
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6288 4146 6316 5528
rect 6366 5400 6422 5409
rect 6472 5370 6500 6734
rect 6564 6361 6592 12038
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6656 9926 6684 11630
rect 6932 10713 6960 14311
rect 7380 14282 7432 14288
rect 7010 13424 7066 13433
rect 7010 13359 7066 13368
rect 7024 13326 7052 13359
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7208 12238 7236 12718
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7116 11830 7144 12106
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7116 11257 7144 11766
rect 7102 11248 7158 11257
rect 7102 11183 7158 11192
rect 7194 11112 7250 11121
rect 7194 11047 7196 11056
rect 7248 11047 7250 11056
rect 7196 11018 7248 11024
rect 7010 10976 7066 10985
rect 7010 10911 7066 10920
rect 6918 10704 6974 10713
rect 6918 10639 6974 10648
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6642 6760 6698 6769
rect 6642 6695 6698 6704
rect 6550 6352 6606 6361
rect 6550 6287 6606 6296
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6366 5335 6422 5344
rect 6460 5364 6512 5370
rect 6092 4140 6144 4146
rect 6276 4140 6328 4146
rect 6092 4082 6144 4088
rect 6196 4100 6276 4128
rect 5446 3703 5502 3712
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 6104 3641 6132 4082
rect 6090 3632 6146 3641
rect 6196 3602 6224 4100
rect 6276 4082 6328 4088
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6090 3567 6146 3576
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 5538 3360 5594 3369
rect 5538 3295 5594 3304
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5354 3088 5410 3097
rect 5172 3052 5224 3058
rect 5354 3023 5356 3032
rect 5172 2994 5224 3000
rect 5408 3023 5410 3032
rect 5356 2994 5408 3000
rect 5552 2938 5580 3295
rect 6090 3224 6146 3233
rect 6090 3159 6146 3168
rect 5460 2910 5580 2938
rect 5460 2530 5488 2910
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5368 2502 5488 2530
rect 5552 2514 5580 2790
rect 5906 2680 5962 2689
rect 5906 2615 5962 2624
rect 5632 2576 5684 2582
rect 5630 2544 5632 2553
rect 5684 2544 5686 2553
rect 5540 2508 5592 2514
rect 5368 2106 5396 2502
rect 5630 2479 5686 2488
rect 5540 2450 5592 2456
rect 5920 2446 5948 2615
rect 5908 2440 5960 2446
rect 5446 2408 5502 2417
rect 5908 2382 5960 2388
rect 5446 2343 5502 2352
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 5460 1970 5488 2343
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 5644 2009 5672 2042
rect 5630 2000 5686 2009
rect 5448 1964 5500 1970
rect 5630 1935 5686 1944
rect 5448 1906 5500 1912
rect 6012 1737 6040 2246
rect 6104 1970 6132 3159
rect 6196 2774 6224 3538
rect 6288 3194 6316 3946
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6380 3058 6408 5335
rect 6460 5306 6512 5312
rect 6564 5302 6592 5782
rect 6552 5296 6604 5302
rect 6472 5244 6552 5250
rect 6472 5238 6604 5244
rect 6472 5222 6592 5238
rect 6472 4214 6500 5222
rect 6656 5114 6684 6695
rect 6748 5302 6776 10474
rect 7024 9994 7052 10911
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7102 10160 7158 10169
rect 7102 10095 7158 10104
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6828 9920 6880 9926
rect 6880 9868 6960 9874
rect 6828 9862 6960 9868
rect 6840 9846 6960 9862
rect 6932 8498 6960 9846
rect 7116 9042 7144 10095
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7116 8362 7144 8978
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6840 5352 6868 6190
rect 6932 5914 6960 7278
rect 7024 6322 7052 7686
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7116 7177 7144 7414
rect 7102 7168 7158 7177
rect 7102 7103 7158 7112
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6920 5364 6972 5370
rect 6840 5324 6920 5352
rect 6920 5306 6972 5312
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6564 5086 6684 5114
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6564 4146 6592 5086
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6656 3126 6684 4966
rect 6840 4622 6868 5102
rect 6828 4616 6880 4622
rect 6734 4584 6790 4593
rect 6828 4558 6880 4564
rect 6734 4519 6790 4528
rect 6748 4486 6776 4519
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 7116 4282 7144 6666
rect 7208 6089 7236 10678
rect 7392 9654 7420 14282
rect 7566 13628 7874 13637
rect 7566 13626 7572 13628
rect 7628 13626 7652 13628
rect 7708 13626 7732 13628
rect 7788 13626 7812 13628
rect 7868 13626 7874 13628
rect 7628 13574 7630 13626
rect 7810 13574 7812 13626
rect 7566 13572 7572 13574
rect 7628 13572 7652 13574
rect 7708 13572 7732 13574
rect 7788 13572 7812 13574
rect 7868 13572 7874 13574
rect 7566 13563 7874 13572
rect 7470 13288 7526 13297
rect 7470 13223 7526 13232
rect 7484 11082 7512 13223
rect 7944 13161 7972 15014
rect 8114 14784 8170 14793
rect 8114 14719 8170 14728
rect 8128 14006 8156 14719
rect 8220 14414 8248 15030
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8404 14482 8432 14894
rect 8956 14521 8984 14962
rect 8942 14512 8998 14521
rect 8392 14476 8444 14482
rect 8942 14447 8998 14456
rect 8392 14418 8444 14424
rect 8208 14408 8260 14414
rect 8260 14368 8340 14396
rect 8208 14350 8260 14356
rect 8206 14104 8262 14113
rect 8206 14039 8262 14048
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 8024 13728 8076 13734
rect 8220 13705 8248 14039
rect 8024 13670 8076 13676
rect 8206 13696 8262 13705
rect 7930 13152 7986 13161
rect 7930 13087 7986 13096
rect 7944 12850 7972 13087
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7944 12646 7972 12786
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7566 12540 7874 12549
rect 7566 12538 7572 12540
rect 7628 12538 7652 12540
rect 7708 12538 7732 12540
rect 7788 12538 7812 12540
rect 7868 12538 7874 12540
rect 7628 12486 7630 12538
rect 7810 12486 7812 12538
rect 7566 12484 7572 12486
rect 7628 12484 7652 12486
rect 7708 12484 7732 12486
rect 7788 12484 7812 12486
rect 7868 12484 7874 12486
rect 7566 12475 7874 12484
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7576 11898 7604 12174
rect 7944 12170 7972 12582
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7566 11452 7874 11461
rect 7566 11450 7572 11452
rect 7628 11450 7652 11452
rect 7708 11450 7732 11452
rect 7788 11450 7812 11452
rect 7868 11450 7874 11452
rect 7628 11398 7630 11450
rect 7810 11398 7812 11450
rect 7566 11396 7572 11398
rect 7628 11396 7652 11398
rect 7708 11396 7732 11398
rect 7788 11396 7812 11398
rect 7868 11396 7874 11398
rect 7566 11387 7874 11396
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7194 6080 7250 6089
rect 7194 6015 7250 6024
rect 7300 4865 7328 8910
rect 7392 7886 7420 9590
rect 7484 7993 7512 11018
rect 8036 10554 8064 13670
rect 8206 13631 8262 13640
rect 8312 12986 8340 14368
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8496 13938 8524 14214
rect 8566 14172 8874 14181
rect 8566 14170 8572 14172
rect 8628 14170 8652 14172
rect 8708 14170 8732 14172
rect 8788 14170 8812 14172
rect 8868 14170 8874 14172
rect 8628 14118 8630 14170
rect 8810 14118 8812 14170
rect 8566 14116 8572 14118
rect 8628 14116 8652 14118
rect 8708 14116 8732 14118
rect 8788 14116 8812 14118
rect 8868 14116 8874 14118
rect 8566 14107 8874 14116
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 8944 13864 8996 13870
rect 8942 13832 8944 13841
rect 8996 13832 8998 13841
rect 8942 13767 8998 13776
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8206 12880 8262 12889
rect 8206 12815 8262 12824
rect 8220 12617 8248 12815
rect 8206 12608 8262 12617
rect 8206 12543 8262 12552
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8220 11082 8248 12106
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8312 10674 8340 12038
rect 8404 10849 8432 13262
rect 8566 13084 8874 13093
rect 8566 13082 8572 13084
rect 8628 13082 8652 13084
rect 8708 13082 8732 13084
rect 8788 13082 8812 13084
rect 8868 13082 8874 13084
rect 8628 13030 8630 13082
rect 8810 13030 8812 13082
rect 8566 13028 8572 13030
rect 8628 13028 8652 13030
rect 8708 13028 8732 13030
rect 8788 13028 8812 13030
rect 8868 13028 8874 13030
rect 8566 13019 8874 13028
rect 8758 12336 8814 12345
rect 8758 12271 8814 12280
rect 8772 12238 8800 12271
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8566 11996 8874 12005
rect 8566 11994 8572 11996
rect 8628 11994 8652 11996
rect 8708 11994 8732 11996
rect 8788 11994 8812 11996
rect 8868 11994 8874 11996
rect 8628 11942 8630 11994
rect 8810 11942 8812 11994
rect 8566 11940 8572 11942
rect 8628 11940 8652 11942
rect 8708 11940 8732 11942
rect 8788 11940 8812 11942
rect 8868 11940 8874 11942
rect 8566 11931 8874 11940
rect 9048 11898 9076 15438
rect 11058 15399 11114 15408
rect 9128 15360 9180 15366
rect 9126 15328 9128 15337
rect 9180 15328 9182 15337
rect 9126 15263 9182 15272
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9140 14385 9168 14758
rect 9220 14408 9272 14414
rect 9126 14376 9182 14385
rect 9220 14350 9272 14356
rect 9126 14311 9182 14320
rect 9126 14104 9182 14113
rect 9126 14039 9128 14048
rect 9180 14039 9182 14048
rect 9128 14010 9180 14016
rect 9232 13025 9260 14350
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9312 14272 9364 14278
rect 9310 14240 9312 14249
rect 9364 14240 9366 14249
rect 9310 14175 9366 14184
rect 9218 13016 9274 13025
rect 9218 12951 9274 12960
rect 9416 12170 9444 14282
rect 11072 14113 11100 15399
rect 12346 14512 12402 14521
rect 12346 14447 12402 14456
rect 10782 14104 10838 14113
rect 10782 14039 10838 14048
rect 11058 14104 11114 14113
rect 11058 14039 11114 14048
rect 9678 13560 9734 13569
rect 9678 13495 9734 13504
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9034 11792 9090 11801
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8944 11756 8996 11762
rect 9034 11727 9090 11736
rect 8944 11698 8996 11704
rect 8772 11529 8800 11698
rect 8758 11520 8814 11529
rect 8758 11455 8814 11464
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8390 10840 8446 10849
rect 8390 10775 8446 10784
rect 8390 10704 8446 10713
rect 8300 10668 8352 10674
rect 8390 10639 8392 10648
rect 8300 10610 8352 10616
rect 8444 10639 8446 10648
rect 8392 10610 8444 10616
rect 8036 10526 8340 10554
rect 7566 10364 7874 10373
rect 7566 10362 7572 10364
rect 7628 10362 7652 10364
rect 7708 10362 7732 10364
rect 7788 10362 7812 10364
rect 7868 10362 7874 10364
rect 7628 10310 7630 10362
rect 7810 10310 7812 10362
rect 7566 10308 7572 10310
rect 7628 10308 7652 10310
rect 7708 10308 7732 10310
rect 7788 10308 7812 10310
rect 7868 10308 7874 10310
rect 7566 10299 7874 10308
rect 8116 10056 8168 10062
rect 8022 10024 8078 10033
rect 8116 9998 8168 10004
rect 8022 9959 8078 9968
rect 8036 9926 8064 9959
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7566 9276 7874 9285
rect 7566 9274 7572 9276
rect 7628 9274 7652 9276
rect 7708 9274 7732 9276
rect 7788 9274 7812 9276
rect 7868 9274 7874 9276
rect 7628 9222 7630 9274
rect 7810 9222 7812 9274
rect 7566 9220 7572 9222
rect 7628 9220 7652 9222
rect 7708 9220 7732 9222
rect 7788 9220 7812 9222
rect 7868 9220 7874 9222
rect 7566 9211 7874 9220
rect 7566 8188 7874 8197
rect 7566 8186 7572 8188
rect 7628 8186 7652 8188
rect 7708 8186 7732 8188
rect 7788 8186 7812 8188
rect 7868 8186 7874 8188
rect 7628 8134 7630 8186
rect 7810 8134 7812 8186
rect 7566 8132 7572 8134
rect 7628 8132 7652 8134
rect 7708 8132 7732 8134
rect 7788 8132 7812 8134
rect 7868 8132 7874 8134
rect 7566 8123 7874 8132
rect 7470 7984 7526 7993
rect 7470 7919 7526 7928
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8036 7546 8064 7822
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7566 7100 7874 7109
rect 7566 7098 7572 7100
rect 7628 7098 7652 7100
rect 7708 7098 7732 7100
rect 7788 7098 7812 7100
rect 7868 7098 7874 7100
rect 7628 7046 7630 7098
rect 7810 7046 7812 7098
rect 7566 7044 7572 7046
rect 7628 7044 7652 7046
rect 7708 7044 7732 7046
rect 7788 7044 7812 7046
rect 7868 7044 7874 7046
rect 7566 7035 7874 7044
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7286 4856 7342 4865
rect 7392 4826 7420 6326
rect 7286 4791 7342 4800
rect 7380 4820 7432 4826
rect 7300 4604 7328 4791
rect 7380 4762 7432 4768
rect 7380 4616 7432 4622
rect 7300 4576 7380 4604
rect 7380 4558 7432 4564
rect 7286 4448 7342 4457
rect 7286 4383 7342 4392
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7010 3632 7066 3641
rect 7010 3567 7066 3576
rect 7024 3534 7052 3567
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7194 3496 7250 3505
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6564 2990 6592 3021
rect 6552 2984 6604 2990
rect 6550 2952 6552 2961
rect 6604 2952 6606 2961
rect 6550 2887 6606 2896
rect 6196 2746 6316 2774
rect 6288 2446 6316 2746
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 6288 1970 6316 2382
rect 6092 1964 6144 1970
rect 6092 1906 6144 1912
rect 6276 1964 6328 1970
rect 6276 1906 6328 1912
rect 6184 1760 6236 1766
rect 5998 1728 6054 1737
rect 6184 1702 6236 1708
rect 5998 1663 6054 1672
rect 6196 1465 6224 1702
rect 6182 1456 6238 1465
rect 6182 1391 6238 1400
rect 6288 1358 6316 1906
rect 6564 1562 6592 2887
rect 6642 2544 6698 2553
rect 6642 2479 6698 2488
rect 6656 2106 6684 2479
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6748 2145 6776 2246
rect 6734 2136 6790 2145
rect 6644 2100 6696 2106
rect 6734 2071 6790 2080
rect 6644 2042 6696 2048
rect 6840 1970 6868 2246
rect 6828 1964 6880 1970
rect 6932 1952 6960 3470
rect 7194 3431 7250 3440
rect 7208 3398 7236 3431
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7300 2774 7328 4383
rect 7392 4282 7420 4558
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7484 3194 7512 6734
rect 7566 6012 7874 6021
rect 7566 6010 7572 6012
rect 7628 6010 7652 6012
rect 7708 6010 7732 6012
rect 7788 6010 7812 6012
rect 7868 6010 7874 6012
rect 7628 5958 7630 6010
rect 7810 5958 7812 6010
rect 7566 5956 7572 5958
rect 7628 5956 7652 5958
rect 7708 5956 7732 5958
rect 7788 5956 7812 5958
rect 7868 5956 7874 5958
rect 7566 5947 7874 5956
rect 7746 5808 7802 5817
rect 7746 5743 7802 5752
rect 7760 5710 7788 5743
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 7566 4924 7874 4933
rect 7566 4922 7572 4924
rect 7628 4922 7652 4924
rect 7708 4922 7732 4924
rect 7788 4922 7812 4924
rect 7868 4922 7874 4924
rect 7628 4870 7630 4922
rect 7810 4870 7812 4922
rect 7566 4868 7572 4870
rect 7628 4868 7652 4870
rect 7708 4868 7732 4870
rect 7788 4868 7812 4870
rect 7868 4868 7874 4870
rect 7566 4859 7874 4868
rect 7566 3836 7874 3845
rect 7566 3834 7572 3836
rect 7628 3834 7652 3836
rect 7708 3834 7732 3836
rect 7788 3834 7812 3836
rect 7868 3834 7874 3836
rect 7628 3782 7630 3834
rect 7810 3782 7812 3834
rect 7566 3780 7572 3782
rect 7628 3780 7652 3782
rect 7708 3780 7732 3782
rect 7788 3780 7812 3782
rect 7868 3780 7874 3782
rect 7566 3771 7874 3780
rect 7944 3618 7972 5578
rect 7852 3590 7972 3618
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7852 2922 7880 3590
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7944 3369 7972 3402
rect 7930 3360 7986 3369
rect 7930 3295 7986 3304
rect 8036 3194 8064 7346
rect 8128 6914 8156 9998
rect 8312 9926 8340 10526
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8298 9752 8354 9761
rect 8298 9687 8354 9696
rect 8206 9208 8262 9217
rect 8206 9143 8262 9152
rect 8220 8430 8248 9143
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8128 6886 8248 6914
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8128 5953 8156 6054
rect 8114 5944 8170 5953
rect 8114 5879 8170 5888
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8128 4690 8156 5714
rect 8220 5522 8248 6886
rect 8312 5914 8340 9687
rect 8404 7313 8432 10610
rect 8496 9625 8524 11086
rect 8566 10908 8874 10917
rect 8566 10906 8572 10908
rect 8628 10906 8652 10908
rect 8708 10906 8732 10908
rect 8788 10906 8812 10908
rect 8868 10906 8874 10908
rect 8628 10854 8630 10906
rect 8810 10854 8812 10906
rect 8566 10852 8572 10854
rect 8628 10852 8652 10854
rect 8708 10852 8732 10854
rect 8788 10852 8812 10854
rect 8868 10852 8874 10854
rect 8566 10843 8874 10852
rect 8956 10266 8984 11698
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8566 9820 8874 9829
rect 8566 9818 8572 9820
rect 8628 9818 8652 9820
rect 8708 9818 8732 9820
rect 8788 9818 8812 9820
rect 8868 9818 8874 9820
rect 8628 9766 8630 9818
rect 8810 9766 8812 9818
rect 8566 9764 8572 9766
rect 8628 9764 8652 9766
rect 8708 9764 8732 9766
rect 8788 9764 8812 9766
rect 8868 9764 8874 9766
rect 8566 9755 8874 9764
rect 8482 9616 8538 9625
rect 8482 9551 8538 9560
rect 9048 9466 9076 11727
rect 9324 11393 9352 12038
rect 9310 11384 9366 11393
rect 9310 11319 9366 11328
rect 9126 10704 9182 10713
rect 9126 10639 9182 10648
rect 9140 10266 9168 10639
rect 9508 10441 9536 12582
rect 9494 10432 9550 10441
rect 9494 10367 9550 10376
rect 9692 10282 9720 13495
rect 10322 13152 10378 13161
rect 10322 13087 10378 13096
rect 9862 11656 9918 11665
rect 9862 11591 9918 11600
rect 9876 10985 9904 11591
rect 10336 11121 10364 13087
rect 10322 11112 10378 11121
rect 10322 11047 10378 11056
rect 9862 10976 9918 10985
rect 9862 10911 9918 10920
rect 10506 10704 10562 10713
rect 10506 10639 10562 10648
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9508 10254 9720 10282
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9324 9722 9352 9930
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 8956 9438 9076 9466
rect 8566 8732 8874 8741
rect 8566 8730 8572 8732
rect 8628 8730 8652 8732
rect 8708 8730 8732 8732
rect 8788 8730 8812 8732
rect 8868 8730 8874 8732
rect 8628 8678 8630 8730
rect 8810 8678 8812 8730
rect 8566 8676 8572 8678
rect 8628 8676 8652 8678
rect 8708 8676 8732 8678
rect 8788 8676 8812 8678
rect 8868 8676 8874 8678
rect 8566 8667 8874 8676
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8390 7304 8446 7313
rect 8390 7239 8446 7248
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8404 5710 8432 7239
rect 8496 6769 8524 7822
rect 8566 7644 8874 7653
rect 8566 7642 8572 7644
rect 8628 7642 8652 7644
rect 8708 7642 8732 7644
rect 8788 7642 8812 7644
rect 8868 7642 8874 7644
rect 8628 7590 8630 7642
rect 8810 7590 8812 7642
rect 8566 7588 8572 7590
rect 8628 7588 8652 7590
rect 8708 7588 8732 7590
rect 8788 7588 8812 7590
rect 8868 7588 8874 7590
rect 8566 7579 8874 7588
rect 8956 7290 8984 9438
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 8974 9076 9318
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9140 8566 9168 8774
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 9126 8392 9182 8401
rect 9126 8327 9182 8336
rect 9140 7546 9168 8327
rect 9508 7886 9536 10254
rect 10520 10130 10548 10639
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8956 7262 9076 7290
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8482 6760 8538 6769
rect 8482 6695 8538 6704
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8220 5494 8340 5522
rect 8206 5400 8262 5409
rect 8206 5335 8208 5344
rect 8260 5335 8262 5344
rect 8208 5306 8260 5312
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8220 4457 8248 5170
rect 8312 4826 8340 5494
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8206 4448 8262 4457
rect 8206 4383 8262 4392
rect 8496 4146 8524 6598
rect 8566 6556 8874 6565
rect 8566 6554 8572 6556
rect 8628 6554 8652 6556
rect 8708 6554 8732 6556
rect 8788 6554 8812 6556
rect 8868 6554 8874 6556
rect 8628 6502 8630 6554
rect 8810 6502 8812 6554
rect 8566 6500 8572 6502
rect 8628 6500 8652 6502
rect 8708 6500 8732 6502
rect 8788 6500 8812 6502
rect 8868 6500 8874 6502
rect 8566 6491 8874 6500
rect 8850 6352 8906 6361
rect 8850 6287 8906 6296
rect 8864 5642 8892 6287
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8566 5468 8874 5477
rect 8566 5466 8572 5468
rect 8628 5466 8652 5468
rect 8708 5466 8732 5468
rect 8788 5466 8812 5468
rect 8868 5466 8874 5468
rect 8628 5414 8630 5466
rect 8810 5414 8812 5466
rect 8566 5412 8572 5414
rect 8628 5412 8652 5414
rect 8708 5412 8732 5414
rect 8788 5412 8812 5414
rect 8868 5412 8874 5414
rect 8566 5403 8874 5412
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 8588 4622 8616 5238
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8566 4380 8874 4389
rect 8566 4378 8572 4380
rect 8628 4378 8652 4380
rect 8708 4378 8732 4380
rect 8788 4378 8812 4380
rect 8868 4378 8874 4380
rect 8628 4326 8630 4378
rect 8810 4326 8812 4378
rect 8566 4324 8572 4326
rect 8628 4324 8652 4326
rect 8708 4324 8732 4326
rect 8788 4324 8812 4326
rect 8868 4324 8874 4326
rect 8566 4315 8874 4324
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8206 3768 8262 3777
rect 8206 3703 8262 3712
rect 8220 3534 8248 3703
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 7208 2746 7328 2774
rect 7566 2748 7874 2757
rect 7566 2746 7572 2748
rect 7628 2746 7652 2748
rect 7708 2746 7732 2748
rect 7788 2746 7812 2748
rect 7868 2746 7874 2748
rect 7208 2446 7236 2746
rect 7628 2694 7630 2746
rect 7810 2694 7812 2746
rect 7566 2692 7572 2694
rect 7628 2692 7652 2694
rect 7708 2692 7732 2694
rect 7788 2692 7812 2694
rect 7868 2692 7874 2694
rect 7566 2683 7874 2692
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 8128 2038 8156 3334
rect 8312 3233 8340 3538
rect 8956 3534 8984 7142
rect 9048 6798 9076 7262
rect 9232 6798 9260 7754
rect 9310 7440 9366 7449
rect 9310 7375 9312 7384
rect 9364 7375 9366 7384
rect 9312 7346 9364 7352
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9048 5778 9076 6734
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8566 3292 8874 3301
rect 8566 3290 8572 3292
rect 8628 3290 8652 3292
rect 8708 3290 8732 3292
rect 8788 3290 8812 3292
rect 8868 3290 8874 3292
rect 8628 3238 8630 3290
rect 8810 3238 8812 3290
rect 8566 3236 8572 3238
rect 8628 3236 8652 3238
rect 8708 3236 8732 3238
rect 8788 3236 8812 3238
rect 8868 3236 8874 3238
rect 8298 3224 8354 3233
rect 8566 3227 8874 3236
rect 8298 3159 8354 3168
rect 9048 3058 9076 5510
rect 9140 4729 9168 6054
rect 9232 5846 9260 6734
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9232 5302 9260 5646
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9126 4720 9182 4729
rect 9126 4655 9182 4664
rect 9220 3936 9272 3942
rect 9218 3904 9220 3913
rect 9272 3904 9274 3913
rect 9218 3839 9274 3848
rect 9218 3496 9274 3505
rect 9218 3431 9274 3440
rect 9232 3398 9260 3431
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9126 3224 9182 3233
rect 9126 3159 9182 3168
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 9034 2952 9090 2961
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8220 2446 8248 2790
rect 8588 2650 8616 2926
rect 9140 2938 9168 3159
rect 9090 2910 9168 2938
rect 9218 2952 9274 2961
rect 9034 2887 9090 2896
rect 9218 2887 9220 2896
rect 9272 2887 9274 2896
rect 9220 2858 9272 2864
rect 8758 2816 8814 2825
rect 8758 2751 8814 2760
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8208 2440 8260 2446
rect 8772 2417 8800 2751
rect 9218 2680 9274 2689
rect 9218 2615 9274 2624
rect 9128 2440 9180 2446
rect 8208 2382 8260 2388
rect 8758 2408 8814 2417
rect 8300 2372 8352 2378
rect 8758 2343 8814 2352
rect 8942 2408 8998 2417
rect 9128 2382 9180 2388
rect 8942 2343 8998 2352
rect 8300 2314 8352 2320
rect 8116 2032 8168 2038
rect 8116 1974 8168 1980
rect 7012 1964 7064 1970
rect 6932 1924 7012 1952
rect 6828 1906 6880 1912
rect 7012 1906 7064 1912
rect 7470 1864 7526 1873
rect 7470 1799 7472 1808
rect 7524 1799 7526 1808
rect 7472 1770 7524 1776
rect 7566 1660 7874 1669
rect 7566 1658 7572 1660
rect 7628 1658 7652 1660
rect 7708 1658 7732 1660
rect 7788 1658 7812 1660
rect 7868 1658 7874 1660
rect 7628 1606 7630 1658
rect 7810 1606 7812 1658
rect 7566 1604 7572 1606
rect 7628 1604 7652 1606
rect 7708 1604 7732 1606
rect 7788 1604 7812 1606
rect 7868 1604 7874 1606
rect 7566 1595 7874 1604
rect 6552 1556 6604 1562
rect 6552 1498 6604 1504
rect 3608 1352 3660 1358
rect 3606 1320 3608 1329
rect 4160 1352 4212 1358
rect 3660 1320 3662 1329
rect 3240 1284 3292 1290
rect 3606 1255 3662 1264
rect 4066 1320 4122 1329
rect 4160 1294 4212 1300
rect 5080 1352 5132 1358
rect 5080 1294 5132 1300
rect 6276 1352 6328 1358
rect 6276 1294 6328 1300
rect 6736 1352 6788 1358
rect 7380 1352 7432 1358
rect 6736 1294 6788 1300
rect 7378 1320 7380 1329
rect 7432 1320 7434 1329
rect 4066 1255 4068 1264
rect 3240 1226 3292 1232
rect 4120 1255 4122 1264
rect 4068 1226 4120 1232
rect 2870 1184 2926 1193
rect 2870 1119 2926 1128
rect 3566 1116 3874 1125
rect 3566 1114 3572 1116
rect 3628 1114 3652 1116
rect 3708 1114 3732 1116
rect 3788 1114 3812 1116
rect 3868 1114 3874 1116
rect 3628 1062 3630 1114
rect 3810 1062 3812 1114
rect 3566 1060 3572 1062
rect 3628 1060 3652 1062
rect 3708 1060 3732 1062
rect 3788 1060 3812 1062
rect 3868 1060 3874 1062
rect 3566 1051 3874 1060
rect 1030 912 1086 921
rect 1030 847 1086 856
rect 4172 649 4200 1294
rect 4344 1216 4396 1222
rect 4344 1158 4396 1164
rect 4896 1216 4948 1222
rect 4896 1158 4948 1164
rect 6000 1216 6052 1222
rect 6000 1158 6052 1164
rect 4356 785 4384 1158
rect 4908 921 4936 1158
rect 6012 1057 6040 1158
rect 5998 1048 6054 1057
rect 5998 983 6054 992
rect 4894 912 4950 921
rect 4894 847 4950 856
rect 4342 776 4398 785
rect 4342 711 4398 720
rect 4158 640 4214 649
rect 4158 575 4214 584
rect 6748 377 6776 1294
rect 7378 1255 7434 1264
rect 8206 1320 8262 1329
rect 8206 1255 8208 1264
rect 8260 1255 8262 1264
rect 8208 1226 8260 1232
rect 8312 649 8340 2314
rect 8390 2272 8446 2281
rect 8390 2207 8446 2216
rect 8404 1737 8432 2207
rect 8566 2204 8874 2213
rect 8566 2202 8572 2204
rect 8628 2202 8652 2204
rect 8708 2202 8732 2204
rect 8788 2202 8812 2204
rect 8868 2202 8874 2204
rect 8628 2150 8630 2202
rect 8810 2150 8812 2202
rect 8566 2148 8572 2150
rect 8628 2148 8652 2150
rect 8708 2148 8732 2150
rect 8788 2148 8812 2150
rect 8868 2148 8874 2150
rect 8566 2139 8874 2148
rect 8956 2106 8984 2343
rect 9034 2272 9090 2281
rect 9034 2207 9090 2216
rect 8944 2100 8996 2106
rect 8944 2042 8996 2048
rect 9048 1970 9076 2207
rect 9036 1964 9088 1970
rect 9036 1906 9088 1912
rect 8390 1728 8446 1737
rect 8390 1663 8446 1672
rect 8566 1116 8874 1125
rect 8566 1114 8572 1116
rect 8628 1114 8652 1116
rect 8708 1114 8732 1116
rect 8788 1114 8812 1116
rect 8868 1114 8874 1116
rect 8628 1062 8630 1114
rect 8810 1062 8812 1114
rect 8566 1060 8572 1062
rect 8628 1060 8652 1062
rect 8708 1060 8732 1062
rect 8788 1060 8812 1062
rect 8868 1060 8874 1062
rect 8566 1051 8874 1060
rect 8114 640 8170 649
rect 8114 575 8170 584
rect 8298 640 8354 649
rect 8298 575 8354 584
rect 6734 368 6790 377
rect 6734 303 6790 312
rect 8128 241 8156 575
rect 9140 513 9168 2382
rect 9232 2106 9260 2615
rect 9324 2446 9352 6598
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9402 5536 9458 5545
rect 9402 5471 9458 5480
rect 9416 4826 9444 5471
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9508 2774 9536 6258
rect 9416 2746 9536 2774
rect 9416 2650 9444 2746
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9600 2145 9628 8366
rect 9692 4622 9720 10066
rect 9770 9072 9826 9081
rect 9770 9007 9826 9016
rect 9784 5234 9812 9007
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9770 4992 9826 5001
rect 9770 4927 9826 4936
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9784 3641 9812 4927
rect 9770 3632 9826 3641
rect 9770 3567 9826 3576
rect 9876 3194 9904 7686
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 9954 5400 10010 5409
rect 9954 5335 9956 5344
rect 10008 5335 10010 5344
rect 9956 5306 10008 5312
rect 9954 3632 10010 3641
rect 9954 3567 9956 3576
rect 10008 3567 10010 3576
rect 9956 3538 10008 3544
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10060 3126 10088 5578
rect 10796 4010 10824 14039
rect 11058 13832 11114 13841
rect 11058 13767 11114 13776
rect 10966 8256 11022 8265
rect 10966 8191 11022 8200
rect 10980 5953 11008 8191
rect 10966 5944 11022 5953
rect 10966 5879 11022 5888
rect 11072 5681 11100 13767
rect 12360 13297 12388 14447
rect 12806 14240 12862 14249
rect 12806 14175 12808 14184
rect 12860 14175 12862 14184
rect 12808 14146 12860 14152
rect 12438 13968 12494 13977
rect 12438 13903 12494 13912
rect 12346 13288 12402 13297
rect 12346 13223 12402 13232
rect 12346 12880 12402 12889
rect 12346 12815 12402 12824
rect 12360 12238 12388 12815
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11150 6488 11206 6497
rect 11150 6423 11206 6432
rect 11058 5672 11114 5681
rect 11058 5607 11114 5616
rect 11164 5273 11192 6423
rect 11150 5264 11206 5273
rect 11150 5199 11206 5208
rect 11058 5128 11114 5137
rect 11058 5063 11114 5072
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10888 2961 10916 4218
rect 11072 3369 11100 5063
rect 11058 3360 11114 3369
rect 11058 3295 11114 3304
rect 10874 2952 10930 2961
rect 10874 2887 10930 2896
rect 9310 2136 9366 2145
rect 9220 2100 9272 2106
rect 9310 2071 9366 2080
rect 9586 2136 9642 2145
rect 9586 2071 9642 2080
rect 9220 2042 9272 2048
rect 9324 1970 9352 2071
rect 9312 1964 9364 1970
rect 9312 1906 9364 1912
rect 11256 1873 11284 8434
rect 11702 7848 11758 7857
rect 11702 7783 11758 7792
rect 11336 7676 11388 7682
rect 11336 7618 11388 7624
rect 11348 5817 11376 7618
rect 11518 6624 11574 6633
rect 11518 6559 11574 6568
rect 11334 5808 11390 5817
rect 11334 5743 11390 5752
rect 11532 3505 11560 6559
rect 11716 5545 11744 7783
rect 11886 7032 11942 7041
rect 11886 6967 11942 6976
rect 11794 6080 11850 6089
rect 11794 6015 11850 6024
rect 11702 5536 11758 5545
rect 11702 5471 11758 5480
rect 11518 3496 11574 3505
rect 11808 3466 11836 6015
rect 11900 4593 11928 6967
rect 12452 6914 12480 13903
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12806 12064 12862 12073
rect 12806 11999 12862 12008
rect 12714 11384 12770 11393
rect 12714 11319 12770 11328
rect 12530 10976 12586 10985
rect 12530 10911 12586 10920
rect 12360 6886 12480 6914
rect 12360 6225 12388 6886
rect 12544 6497 12572 10911
rect 12622 10024 12678 10033
rect 12622 9959 12678 9968
rect 12530 6488 12586 6497
rect 12530 6423 12586 6432
rect 12346 6216 12402 6225
rect 12346 6151 12402 6160
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11886 4584 11942 4593
rect 11886 4519 11942 4528
rect 12070 4584 12126 4593
rect 12070 4519 12126 4528
rect 11518 3431 11574 3440
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11702 3360 11758 3369
rect 11702 3295 11758 3304
rect 11242 1864 11298 1873
rect 11242 1799 11298 1808
rect 11716 1737 11744 3295
rect 12084 2281 12112 4519
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 12268 3233 12296 3402
rect 12254 3224 12310 3233
rect 12254 3159 12310 3168
rect 12360 2825 12388 4762
rect 12636 3777 12664 9959
rect 12728 4865 12756 11319
rect 12714 4856 12770 4865
rect 12714 4791 12770 4800
rect 12622 3768 12678 3777
rect 12622 3703 12678 3712
rect 12820 3641 12848 11999
rect 12898 11520 12954 11529
rect 12898 11455 12954 11464
rect 12806 3632 12862 3641
rect 12806 3567 12862 3576
rect 12912 3466 12940 11455
rect 12900 3460 12952 3466
rect 12900 3402 12952 3408
rect 13004 3369 13032 12174
rect 13096 8974 13124 16079
rect 13450 16008 13506 16017
rect 13634 16008 13690 16017
rect 13450 15943 13506 15952
rect 13556 15966 13634 15994
rect 13464 12889 13492 15943
rect 13450 12880 13506 12889
rect 13450 12815 13506 12824
rect 13450 12744 13506 12753
rect 13450 12679 13452 12688
rect 13504 12679 13506 12688
rect 13452 12650 13504 12656
rect 13556 11830 13584 15966
rect 13634 15943 13690 15952
rect 13634 15328 13690 15337
rect 13634 15263 13636 15272
rect 13688 15263 13690 15272
rect 13636 15234 13688 15240
rect 13634 14920 13690 14929
rect 13634 14855 13636 14864
rect 13688 14855 13690 14864
rect 13636 14826 13688 14832
rect 13634 14784 13690 14793
rect 13634 14719 13636 14728
rect 13688 14719 13690 14728
rect 13636 14690 13688 14696
rect 13634 14648 13690 14657
rect 13634 14583 13636 14592
rect 13688 14583 13690 14592
rect 13636 14554 13688 14560
rect 13740 14385 13768 16623
rect 15120 15178 15148 16623
rect 17912 15600 17968 15609
rect 17968 15558 18092 15586
rect 17912 15535 17968 15544
rect 16488 15292 16540 15298
rect 16488 15234 16540 15240
rect 15120 15150 15240 15178
rect 13820 14816 13872 14822
rect 13818 14784 13820 14793
rect 13872 14784 13874 14793
rect 13818 14719 13874 14728
rect 14188 14748 14240 14754
rect 14188 14690 14240 14696
rect 13726 14376 13782 14385
rect 13726 14311 13782 14320
rect 13634 14240 13690 14249
rect 13634 14175 13690 14184
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 13542 11520 13598 11529
rect 13542 11455 13544 11464
rect 13596 11455 13598 11464
rect 13544 11426 13596 11432
rect 13648 10713 13676 14175
rect 13726 13696 13782 13705
rect 13726 13631 13782 13640
rect 13740 13598 13768 13631
rect 13728 13592 13780 13598
rect 13728 13534 13780 13540
rect 13818 13560 13874 13569
rect 13818 13495 13820 13504
rect 13872 13495 13874 13504
rect 13820 13466 13872 13472
rect 13726 13424 13782 13433
rect 13726 13359 13782 13368
rect 13740 11098 13768 13359
rect 13818 13016 13874 13025
rect 13818 12951 13820 12960
rect 13872 12951 13874 12960
rect 13820 12922 13872 12928
rect 13818 12608 13874 12617
rect 13818 12543 13820 12552
rect 13872 12543 13874 12552
rect 13820 12514 13872 12520
rect 13820 12232 13872 12238
rect 13818 12200 13820 12209
rect 13872 12200 13874 12209
rect 13818 12135 13874 12144
rect 13820 11960 13872 11966
rect 13818 11928 13820 11937
rect 13872 11928 13874 11937
rect 13818 11863 13874 11872
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13832 11257 13860 11766
rect 13818 11248 13874 11257
rect 13818 11183 13874 11192
rect 13740 11070 13860 11098
rect 13634 10704 13690 10713
rect 13634 10639 13690 10648
rect 13542 10568 13598 10577
rect 13832 10538 13860 11070
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 13542 10503 13598 10512
rect 13820 10532 13872 10538
rect 13176 9512 13228 9518
rect 13174 9480 13176 9489
rect 13228 9480 13230 9489
rect 13174 9415 13230 9424
rect 13450 9208 13506 9217
rect 13450 9143 13506 9152
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13280 6089 13308 8230
rect 13266 6080 13322 6089
rect 13266 6015 13322 6024
rect 13464 5001 13492 9143
rect 13556 8362 13584 10503
rect 13820 10474 13872 10480
rect 13818 10432 13874 10441
rect 13874 10390 14044 10418
rect 13818 10367 13874 10376
rect 13820 10328 13872 10334
rect 13818 10296 13820 10305
rect 13872 10296 13874 10305
rect 13818 10231 13874 10240
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13740 9761 13768 10134
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13726 9752 13782 9761
rect 13726 9687 13782 9696
rect 13818 9344 13874 9353
rect 13818 9279 13874 9288
rect 13832 9246 13860 9279
rect 13820 9240 13872 9246
rect 13820 9182 13872 9188
rect 13820 9104 13872 9110
rect 13818 9072 13820 9081
rect 13872 9072 13874 9081
rect 13818 9007 13874 9016
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13820 7472 13872 7478
rect 13818 7440 13820 7449
rect 13872 7440 13874 7449
rect 13818 7375 13874 7384
rect 13818 6896 13874 6905
rect 13818 6831 13874 6840
rect 13832 6798 13860 6831
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13820 5840 13872 5846
rect 13818 5808 13820 5817
rect 13872 5808 13874 5817
rect 13818 5743 13874 5752
rect 13832 5642 13860 5743
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13636 5296 13688 5302
rect 13634 5264 13636 5273
rect 13688 5264 13690 5273
rect 13634 5199 13690 5208
rect 13740 5137 13768 5510
rect 13818 5400 13874 5409
rect 13818 5335 13874 5344
rect 13726 5128 13782 5137
rect 13726 5063 13782 5072
rect 13450 4992 13506 5001
rect 13450 4927 13506 4936
rect 13726 4856 13782 4865
rect 13726 4791 13782 4800
rect 13740 4185 13768 4791
rect 13726 4176 13782 4185
rect 13726 4111 13782 4120
rect 13832 3942 13860 5335
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13818 3768 13874 3777
rect 13818 3703 13874 3712
rect 12990 3360 13046 3369
rect 12990 3295 13046 3304
rect 12346 2816 12402 2825
rect 12346 2751 12402 2760
rect 12070 2272 12126 2281
rect 12070 2207 12126 2216
rect 13832 2009 13860 3703
rect 13818 2000 13874 2009
rect 13818 1935 13874 1944
rect 11702 1728 11758 1737
rect 11702 1663 11758 1672
rect 9126 504 9182 513
rect 9126 439 9182 448
rect 13924 377 13952 9862
rect 14016 2774 14044 10390
rect 14108 9926 14136 10950
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14200 5574 14228 14690
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14844 11082 14872 14554
rect 15212 14414 15240 15150
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15028 12238 15056 12786
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14016 2746 14136 2774
rect 13910 368 13966 377
rect 13910 303 13966 312
rect 14108 241 14136 2746
rect 14292 921 14320 8978
rect 15212 8498 15240 12650
rect 15304 9654 15332 14758
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15396 9042 15424 14418
rect 16028 13592 16080 13598
rect 16028 13534 16080 13540
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15488 11966 15516 13194
rect 15476 11960 15528 11966
rect 15476 11902 15528 11908
rect 15660 11484 15712 11490
rect 15660 11426 15712 11432
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15488 9246 15516 9862
rect 15476 9240 15528 9246
rect 15476 9182 15528 9188
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15396 2774 15424 8842
rect 15580 5846 15608 10066
rect 15672 6798 15700 11426
rect 15764 9110 15792 13398
rect 15936 12572 15988 12578
rect 15936 12514 15988 12520
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15752 9104 15804 9110
rect 15752 9046 15804 9052
rect 15856 7682 15884 12174
rect 15948 8906 15976 12514
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 16040 8294 16068 13534
rect 16500 11830 16528 15234
rect 17912 15192 17968 15201
rect 17912 15127 17914 15136
rect 17966 15127 17968 15136
rect 17914 15098 17966 15104
rect 17408 14884 17460 14890
rect 17408 14826 17460 14832
rect 17132 14204 17184 14210
rect 17132 14146 17184 14152
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 15844 7676 15896 7682
rect 15844 7618 15896 7624
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 15120 2746 15424 2774
rect 15120 1465 15148 2746
rect 16868 2417 16896 3878
rect 16854 2408 16910 2417
rect 16854 2343 16910 2352
rect 16960 1601 16988 10474
rect 17144 5302 17172 14146
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17328 4185 17356 12922
rect 17420 4826 17448 14826
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17314 4176 17370 4185
rect 17314 4111 17370 4120
rect 17604 2786 17632 14350
rect 17914 13592 17966 13598
rect 17912 13560 17914 13569
rect 17966 13560 17968 13569
rect 17912 13495 17968 13504
rect 18064 9518 18092 15558
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17696 5522 17724 8910
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 17912 6216 17968 6225
rect 17912 6151 17914 6160
rect 17966 6151 17968 6160
rect 17914 6122 17966 6128
rect 17696 5494 18000 5522
rect 17972 2938 18000 5494
rect 18064 3913 18092 7414
rect 18050 3904 18106 3913
rect 18050 3839 18106 3848
rect 17972 2910 18092 2938
rect 17592 2780 17644 2786
rect 17592 2722 17644 2728
rect 17960 2780 18012 2786
rect 17960 2722 18012 2728
rect 17972 1714 18000 2722
rect 18064 2553 18092 2910
rect 18050 2544 18106 2553
rect 18050 2479 18106 2488
rect 17788 1686 18000 1714
rect 16946 1592 17002 1601
rect 16946 1527 17002 1536
rect 15106 1456 15162 1465
rect 15106 1391 15162 1400
rect 14278 912 14334 921
rect 14278 847 14334 856
rect 17788 785 17816 1686
rect 18156 1578 18184 11018
rect 18248 4282 18276 16623
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18340 3777 18368 13466
rect 18432 10334 18460 16895
rect 19062 16688 19118 16697
rect 19062 16623 19118 16632
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18420 10328 18472 10334
rect 18420 10270 18472 10276
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18326 3768 18382 3777
rect 18326 3703 18382 3712
rect 18432 2145 18460 10134
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18418 2136 18474 2145
rect 18418 2071 18474 2080
rect 18064 1550 18184 1578
rect 18064 1442 18092 1550
rect 17880 1414 18092 1442
rect 17774 776 17830 785
rect 17774 711 17830 720
rect 17880 649 17908 1414
rect 18524 1329 18552 8298
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18510 1320 18566 1329
rect 18510 1255 18566 1264
rect 17866 640 17922 649
rect 17866 575 17922 584
rect 18616 513 18644 6122
rect 18800 4321 18828 15098
rect 18972 13592 19024 13598
rect 18972 13534 19024 13540
rect 18786 4312 18842 4321
rect 18786 4247 18842 4256
rect 18984 4049 19012 13534
rect 19076 5778 19104 16623
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 19064 5636 19116 5642
rect 19064 5578 19116 5584
rect 18970 4040 19026 4049
rect 18970 3975 19026 3984
rect 19076 3097 19104 5578
rect 19062 3088 19118 3097
rect 19062 3023 19118 3032
rect 18602 504 18658 513
rect 18602 439 18658 448
rect 8114 232 8170 241
rect 8114 167 8170 176
rect 14094 232 14150 241
rect 14094 167 14150 176
<< via2 >>
rect 2410 16904 2466 16960
rect 386 15272 442 15328
rect 202 14456 258 14512
rect 478 14864 534 14920
rect 570 12144 626 12200
rect 294 1536 350 1592
rect 754 9696 810 9752
rect 938 11056 994 11112
rect 1214 13776 1270 13832
rect 1766 15444 1768 15464
rect 1768 15444 1820 15464
rect 1820 15444 1822 15464
rect 1766 15408 1822 15444
rect 3146 16768 3202 16824
rect 2572 15802 2628 15804
rect 2652 15802 2708 15804
rect 2732 15802 2788 15804
rect 2812 15802 2868 15804
rect 2572 15750 2618 15802
rect 2618 15750 2628 15802
rect 2652 15750 2682 15802
rect 2682 15750 2694 15802
rect 2694 15750 2708 15802
rect 2732 15750 2746 15802
rect 2746 15750 2758 15802
rect 2758 15750 2788 15802
rect 2812 15750 2822 15802
rect 2822 15750 2868 15802
rect 2572 15748 2628 15750
rect 2652 15748 2708 15750
rect 2732 15748 2788 15750
rect 2812 15748 2868 15750
rect 2778 15308 2780 15328
rect 2780 15308 2832 15328
rect 2832 15308 2834 15328
rect 2778 15272 2834 15308
rect 1122 9016 1178 9072
rect 1122 8336 1178 8392
rect 1030 7792 1086 7848
rect 938 1400 994 1456
rect 570 1128 626 1184
rect 1306 12008 1362 12064
rect 1582 12416 1638 12472
rect 1398 11600 1454 11656
rect 2226 13232 2282 13288
rect 2134 11736 2190 11792
rect 1582 6840 1638 6896
rect 1398 5208 1454 5264
rect 1306 4664 1362 4720
rect 2778 14884 2834 14920
rect 2778 14864 2780 14884
rect 2780 14864 2832 14884
rect 2832 14864 2834 14884
rect 2572 14714 2628 14716
rect 2652 14714 2708 14716
rect 2732 14714 2788 14716
rect 2812 14714 2868 14716
rect 2572 14662 2618 14714
rect 2618 14662 2628 14714
rect 2652 14662 2682 14714
rect 2682 14662 2694 14714
rect 2694 14662 2708 14714
rect 2732 14662 2746 14714
rect 2746 14662 2758 14714
rect 2758 14662 2788 14714
rect 2812 14662 2822 14714
rect 2822 14662 2868 14714
rect 2572 14660 2628 14662
rect 2652 14660 2708 14662
rect 2732 14660 2788 14662
rect 2812 14660 2868 14662
rect 2502 13912 2558 13968
rect 2778 13776 2834 13832
rect 2572 13626 2628 13628
rect 2652 13626 2708 13628
rect 2732 13626 2788 13628
rect 2812 13626 2868 13628
rect 2572 13574 2618 13626
rect 2618 13574 2628 13626
rect 2652 13574 2682 13626
rect 2682 13574 2694 13626
rect 2694 13574 2708 13626
rect 2732 13574 2746 13626
rect 2746 13574 2758 13626
rect 2758 13574 2788 13626
rect 2812 13574 2822 13626
rect 2822 13574 2868 13626
rect 2572 13572 2628 13574
rect 2652 13572 2708 13574
rect 2732 13572 2788 13574
rect 2812 13572 2868 13574
rect 3146 13912 3202 13968
rect 2594 12724 2596 12744
rect 2596 12724 2648 12744
rect 2648 12724 2650 12744
rect 2594 12688 2650 12724
rect 2572 12538 2628 12540
rect 2652 12538 2708 12540
rect 2732 12538 2788 12540
rect 2812 12538 2868 12540
rect 2572 12486 2618 12538
rect 2618 12486 2628 12538
rect 2652 12486 2682 12538
rect 2682 12486 2694 12538
rect 2694 12486 2708 12538
rect 2732 12486 2746 12538
rect 2746 12486 2758 12538
rect 2758 12486 2788 12538
rect 2812 12486 2822 12538
rect 2822 12486 2868 12538
rect 2572 12484 2628 12486
rect 2652 12484 2708 12486
rect 2732 12484 2788 12486
rect 2812 12484 2868 12486
rect 4710 16632 4766 16688
rect 4066 16088 4122 16144
rect 3572 15258 3628 15260
rect 3652 15258 3708 15260
rect 3732 15258 3788 15260
rect 3812 15258 3868 15260
rect 3572 15206 3618 15258
rect 3618 15206 3628 15258
rect 3652 15206 3682 15258
rect 3682 15206 3694 15258
rect 3694 15206 3708 15258
rect 3732 15206 3746 15258
rect 3746 15206 3758 15258
rect 3758 15206 3788 15258
rect 3812 15206 3822 15258
rect 3822 15206 3868 15258
rect 3572 15204 3628 15206
rect 3652 15204 3708 15206
rect 3732 15204 3788 15206
rect 3812 15204 3868 15206
rect 4066 15020 4122 15056
rect 4066 15000 4068 15020
rect 4068 15000 4120 15020
rect 4120 15000 4122 15020
rect 3974 14356 3976 14376
rect 3976 14356 4028 14376
rect 4028 14356 4030 14376
rect 3974 14320 4030 14356
rect 3572 14170 3628 14172
rect 3652 14170 3708 14172
rect 3732 14170 3788 14172
rect 3812 14170 3868 14172
rect 3572 14118 3618 14170
rect 3618 14118 3628 14170
rect 3652 14118 3682 14170
rect 3682 14118 3694 14170
rect 3694 14118 3708 14170
rect 3732 14118 3746 14170
rect 3746 14118 3758 14170
rect 3758 14118 3788 14170
rect 3812 14118 3822 14170
rect 3822 14118 3868 14170
rect 3572 14116 3628 14118
rect 3652 14116 3708 14118
rect 3732 14116 3788 14118
rect 3812 14116 3868 14118
rect 3422 13368 3478 13424
rect 3572 13082 3628 13084
rect 3652 13082 3708 13084
rect 3732 13082 3788 13084
rect 3812 13082 3868 13084
rect 3572 13030 3618 13082
rect 3618 13030 3628 13082
rect 3652 13030 3682 13082
rect 3682 13030 3694 13082
rect 3694 13030 3708 13082
rect 3732 13030 3746 13082
rect 3746 13030 3758 13082
rect 3758 13030 3788 13082
rect 3812 13030 3822 13082
rect 3822 13030 3868 13082
rect 3572 13028 3628 13030
rect 3652 13028 3708 13030
rect 3732 13028 3788 13030
rect 3812 13028 3868 13030
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2686 11212 2742 11248
rect 2686 11192 2688 11212
rect 2688 11192 2740 11212
rect 2740 11192 2742 11212
rect 2502 10548 2504 10568
rect 2504 10548 2556 10568
rect 2556 10548 2558 10568
rect 2502 10512 2558 10548
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 3514 12144 3570 12200
rect 3572 11994 3628 11996
rect 3652 11994 3708 11996
rect 3732 11994 3788 11996
rect 3812 11994 3868 11996
rect 3572 11942 3618 11994
rect 3618 11942 3628 11994
rect 3652 11942 3682 11994
rect 3682 11942 3694 11994
rect 3694 11942 3708 11994
rect 3732 11942 3746 11994
rect 3746 11942 3758 11994
rect 3758 11942 3788 11994
rect 3812 11942 3822 11994
rect 3822 11942 3868 11994
rect 3572 11940 3628 11942
rect 3652 11940 3708 11942
rect 3732 11940 3788 11942
rect 3812 11940 3868 11942
rect 2962 10104 3018 10160
rect 2686 9460 2688 9480
rect 2688 9460 2740 9480
rect 2740 9460 2742 9480
rect 2686 9424 2742 9460
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2226 7384 2282 7440
rect 2778 8372 2780 8392
rect 2780 8372 2832 8392
rect 2832 8372 2834 8392
rect 2778 8336 2834 8372
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2410 7928 2466 7984
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 3606 11464 3662 11520
rect 3238 11076 3294 11112
rect 3238 11056 3240 11076
rect 3240 11056 3292 11076
rect 3292 11056 3294 11076
rect 3572 10906 3628 10908
rect 3652 10906 3708 10908
rect 3732 10906 3788 10908
rect 3812 10906 3868 10908
rect 3572 10854 3618 10906
rect 3618 10854 3628 10906
rect 3652 10854 3682 10906
rect 3682 10854 3694 10906
rect 3694 10854 3708 10906
rect 3732 10854 3746 10906
rect 3746 10854 3758 10906
rect 3758 10854 3788 10906
rect 3812 10854 3822 10906
rect 3822 10854 3868 10906
rect 3572 10852 3628 10854
rect 3652 10852 3708 10854
rect 3732 10852 3788 10854
rect 3812 10852 3868 10854
rect 3330 9968 3386 10024
rect 3238 9696 3294 9752
rect 3054 7928 3110 7984
rect 3054 6840 3110 6896
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 3238 8880 3294 8936
rect 3238 7248 3294 7304
rect 3054 5888 3110 5944
rect 2502 5652 2504 5672
rect 2504 5652 2556 5672
rect 2556 5652 2558 5672
rect 2502 5616 2558 5652
rect 2410 4800 2466 4856
rect 2410 4120 2466 4176
rect 2410 3984 2466 4040
rect 2686 3984 2742 4040
rect 2594 3848 2650 3904
rect 2686 3712 2742 3768
rect 2502 2624 2558 2680
rect 3146 3848 3202 3904
rect 3146 3576 3202 3632
rect 2686 2488 2742 2544
rect 1858 1536 1914 1592
rect 2318 1536 2374 1592
rect 2870 1672 2926 1728
rect 2778 1400 2834 1456
rect 1122 1264 1178 1320
rect 3572 9818 3628 9820
rect 3652 9818 3708 9820
rect 3732 9818 3788 9820
rect 3812 9818 3868 9820
rect 3572 9766 3618 9818
rect 3618 9766 3628 9818
rect 3652 9766 3682 9818
rect 3682 9766 3694 9818
rect 3694 9766 3708 9818
rect 3732 9766 3746 9818
rect 3746 9766 3758 9818
rect 3758 9766 3788 9818
rect 3812 9766 3822 9818
rect 3822 9766 3868 9818
rect 3572 9764 3628 9766
rect 3652 9764 3708 9766
rect 3732 9764 3788 9766
rect 3812 9764 3868 9766
rect 4066 14184 4122 14240
rect 4066 14048 4122 14104
rect 4066 13096 4122 13152
rect 4158 11636 4160 11656
rect 4160 11636 4212 11656
rect 4212 11636 4214 11656
rect 4158 11600 4214 11636
rect 4066 11056 4122 11112
rect 4434 14492 4436 14512
rect 4436 14492 4488 14512
rect 4488 14492 4490 14512
rect 4434 14456 4490 14492
rect 6182 16224 6238 16280
rect 4434 12960 4490 13016
rect 4342 11872 4398 11928
rect 5262 15408 5318 15464
rect 5722 15952 5778 16008
rect 5354 15000 5410 15056
rect 5446 14864 5502 14920
rect 4894 13932 4950 13968
rect 4894 13912 4896 13932
rect 4896 13912 4948 13932
rect 4948 13912 4950 13932
rect 4342 9968 4398 10024
rect 4066 9152 4122 9208
rect 4526 9696 4582 9752
rect 3572 8730 3628 8732
rect 3652 8730 3708 8732
rect 3732 8730 3788 8732
rect 3812 8730 3868 8732
rect 3572 8678 3618 8730
rect 3618 8678 3628 8730
rect 3652 8678 3682 8730
rect 3682 8678 3694 8730
rect 3694 8678 3708 8730
rect 3732 8678 3746 8730
rect 3746 8678 3758 8730
rect 3758 8678 3788 8730
rect 3812 8678 3822 8730
rect 3822 8678 3868 8730
rect 3572 8676 3628 8678
rect 3652 8676 3708 8678
rect 3732 8676 3788 8678
rect 3812 8676 3868 8678
rect 3882 7948 3938 7984
rect 3882 7928 3884 7948
rect 3884 7928 3936 7948
rect 3936 7928 3938 7948
rect 3514 7792 3570 7848
rect 3572 7642 3628 7644
rect 3652 7642 3708 7644
rect 3732 7642 3788 7644
rect 3812 7642 3868 7644
rect 3572 7590 3618 7642
rect 3618 7590 3628 7642
rect 3652 7590 3682 7642
rect 3682 7590 3694 7642
rect 3694 7590 3708 7642
rect 3732 7590 3746 7642
rect 3746 7590 3758 7642
rect 3758 7590 3788 7642
rect 3812 7590 3822 7642
rect 3822 7590 3868 7642
rect 3572 7588 3628 7590
rect 3652 7588 3708 7590
rect 3732 7588 3788 7590
rect 3812 7588 3868 7590
rect 3572 6554 3628 6556
rect 3652 6554 3708 6556
rect 3732 6554 3788 6556
rect 3812 6554 3868 6556
rect 3572 6502 3618 6554
rect 3618 6502 3628 6554
rect 3652 6502 3682 6554
rect 3682 6502 3694 6554
rect 3694 6502 3708 6554
rect 3732 6502 3746 6554
rect 3746 6502 3758 6554
rect 3758 6502 3788 6554
rect 3812 6502 3822 6554
rect 3822 6502 3868 6554
rect 3572 6500 3628 6502
rect 3652 6500 3708 6502
rect 3732 6500 3788 6502
rect 3812 6500 3868 6502
rect 3514 6296 3570 6352
rect 3572 5466 3628 5468
rect 3652 5466 3708 5468
rect 3732 5466 3788 5468
rect 3812 5466 3868 5468
rect 3572 5414 3618 5466
rect 3618 5414 3628 5466
rect 3652 5414 3682 5466
rect 3682 5414 3694 5466
rect 3694 5414 3708 5466
rect 3732 5414 3746 5466
rect 3746 5414 3758 5466
rect 3758 5414 3788 5466
rect 3812 5414 3822 5466
rect 3822 5414 3868 5466
rect 3572 5412 3628 5414
rect 3652 5412 3708 5414
rect 3732 5412 3788 5414
rect 3812 5412 3868 5414
rect 4066 6976 4122 7032
rect 4158 5072 4214 5128
rect 3514 4664 3570 4720
rect 3572 4378 3628 4380
rect 3652 4378 3708 4380
rect 3732 4378 3788 4380
rect 3812 4378 3868 4380
rect 3572 4326 3618 4378
rect 3618 4326 3628 4378
rect 3652 4326 3682 4378
rect 3682 4326 3694 4378
rect 3694 4326 3708 4378
rect 3732 4326 3746 4378
rect 3746 4326 3758 4378
rect 3758 4326 3788 4378
rect 3812 4326 3822 4378
rect 3822 4326 3868 4378
rect 3572 4324 3628 4326
rect 3652 4324 3708 4326
rect 3732 4324 3788 4326
rect 3812 4324 3868 4326
rect 3974 4120 4030 4176
rect 3330 3848 3386 3904
rect 3572 3290 3628 3292
rect 3652 3290 3708 3292
rect 3732 3290 3788 3292
rect 3812 3290 3868 3292
rect 3572 3238 3618 3290
rect 3618 3238 3628 3290
rect 3652 3238 3682 3290
rect 3682 3238 3694 3290
rect 3694 3238 3708 3290
rect 3732 3238 3746 3290
rect 3746 3238 3758 3290
rect 3758 3238 3788 3290
rect 3812 3238 3822 3290
rect 3822 3238 3868 3290
rect 3572 3236 3628 3238
rect 3652 3236 3708 3238
rect 3732 3236 3788 3238
rect 3812 3236 3868 3238
rect 4066 4020 4068 4040
rect 4068 4020 4120 4040
rect 4120 4020 4122 4040
rect 4066 3984 4122 4020
rect 4342 3848 4398 3904
rect 3572 2202 3628 2204
rect 3652 2202 3708 2204
rect 3732 2202 3788 2204
rect 3812 2202 3868 2204
rect 3572 2150 3618 2202
rect 3618 2150 3628 2202
rect 3652 2150 3682 2202
rect 3682 2150 3694 2202
rect 3694 2150 3708 2202
rect 3732 2150 3746 2202
rect 3746 2150 3758 2202
rect 3758 2150 3788 2202
rect 3812 2150 3822 2202
rect 3822 2150 3868 2202
rect 3572 2148 3628 2150
rect 3652 2148 3708 2150
rect 3732 2148 3788 2150
rect 3812 2148 3868 2150
rect 4526 6704 4582 6760
rect 4894 11464 4950 11520
rect 4802 10804 4858 10840
rect 4802 10784 4804 10804
rect 4804 10784 4856 10804
rect 4856 10784 4858 10804
rect 4986 11056 5042 11112
rect 4986 9016 5042 9072
rect 4618 5888 4674 5944
rect 4618 5752 4674 5808
rect 4526 5208 4582 5264
rect 4802 5616 4858 5672
rect 4986 5616 5042 5672
rect 4710 5208 4766 5264
rect 4710 4664 4766 4720
rect 4894 4800 4950 4856
rect 5538 11736 5594 11792
rect 5446 11192 5502 11248
rect 4158 1536 4214 1592
rect 4710 2252 4712 2272
rect 4712 2252 4764 2272
rect 4764 2252 4766 2272
rect 4710 2216 4766 2252
rect 18418 16904 18474 16960
rect 13634 16768 13690 16824
rect 13726 16632 13782 16688
rect 15106 16632 15162 16688
rect 15290 16668 15292 16688
rect 15292 16668 15344 16688
rect 15344 16668 15346 16688
rect 15290 16632 15346 16668
rect 18234 16632 18290 16688
rect 13082 16088 13138 16144
rect 7572 15802 7628 15804
rect 7652 15802 7708 15804
rect 7732 15802 7788 15804
rect 7812 15802 7868 15804
rect 7572 15750 7618 15802
rect 7618 15750 7628 15802
rect 7652 15750 7682 15802
rect 7682 15750 7694 15802
rect 7694 15750 7708 15802
rect 7732 15750 7746 15802
rect 7746 15750 7758 15802
rect 7758 15750 7788 15802
rect 7812 15750 7822 15802
rect 7822 15750 7868 15802
rect 7572 15748 7628 15750
rect 7652 15748 7708 15750
rect 7732 15748 7788 15750
rect 7812 15748 7868 15750
rect 8114 15428 8170 15464
rect 8114 15408 8116 15428
rect 8116 15408 8168 15428
rect 8168 15408 8170 15428
rect 6550 15136 6606 15192
rect 8572 15258 8628 15260
rect 8652 15258 8708 15260
rect 8732 15258 8788 15260
rect 8812 15258 8868 15260
rect 8572 15206 8618 15258
rect 8618 15206 8628 15258
rect 8652 15206 8682 15258
rect 8682 15206 8694 15258
rect 8694 15206 8708 15258
rect 8732 15206 8746 15258
rect 8746 15206 8758 15258
rect 8758 15206 8788 15258
rect 8812 15206 8822 15258
rect 8822 15206 8868 15258
rect 8572 15204 8628 15206
rect 8652 15204 8708 15206
rect 8732 15204 8788 15206
rect 8812 15204 8868 15206
rect 8390 15136 8446 15192
rect 7572 14714 7628 14716
rect 7652 14714 7708 14716
rect 7732 14714 7788 14716
rect 7812 14714 7868 14716
rect 7572 14662 7618 14714
rect 7618 14662 7628 14714
rect 7652 14662 7682 14714
rect 7682 14662 7694 14714
rect 7694 14662 7708 14714
rect 7732 14662 7746 14714
rect 7746 14662 7758 14714
rect 7758 14662 7788 14714
rect 7812 14662 7822 14714
rect 7822 14662 7868 14714
rect 7572 14660 7628 14662
rect 7652 14660 7708 14662
rect 7732 14660 7788 14662
rect 7812 14660 7868 14662
rect 6918 14320 6974 14376
rect 6642 13812 6644 13832
rect 6644 13812 6696 13832
rect 6696 13812 6698 13832
rect 6642 13776 6698 13812
rect 6642 12824 6698 12880
rect 6090 12280 6146 12336
rect 5998 12144 6054 12200
rect 5630 9696 5686 9752
rect 5630 8472 5686 8528
rect 5354 8336 5410 8392
rect 5354 7112 5410 7168
rect 5446 6024 5502 6080
rect 5446 4936 5502 4992
rect 5446 4800 5502 4856
rect 5262 4256 5318 4312
rect 5814 9560 5870 9616
rect 5814 9152 5870 9208
rect 6274 11600 6330 11656
rect 6366 11464 6422 11520
rect 6090 11328 6146 11384
rect 6458 11056 6514 11112
rect 5998 9696 6054 9752
rect 5998 9288 6054 9344
rect 5998 6160 6054 6216
rect 5906 4256 5962 4312
rect 5446 3712 5502 3768
rect 6366 6976 6422 7032
rect 6274 6432 6330 6488
rect 6182 5752 6238 5808
rect 6182 4664 6238 4720
rect 6366 5344 6422 5400
rect 7010 13368 7066 13424
rect 7102 11192 7158 11248
rect 7194 11076 7250 11112
rect 7194 11056 7196 11076
rect 7196 11056 7248 11076
rect 7248 11056 7250 11076
rect 7010 10920 7066 10976
rect 6918 10648 6974 10704
rect 6642 6704 6698 6760
rect 6550 6296 6606 6352
rect 6090 3576 6146 3632
rect 5538 3304 5594 3360
rect 5354 3052 5410 3088
rect 5354 3032 5356 3052
rect 5356 3032 5408 3052
rect 5408 3032 5410 3052
rect 6090 3168 6146 3224
rect 5906 2624 5962 2680
rect 5630 2524 5632 2544
rect 5632 2524 5684 2544
rect 5684 2524 5686 2544
rect 5630 2488 5686 2524
rect 5446 2352 5502 2408
rect 5630 1944 5686 2000
rect 7102 10104 7158 10160
rect 7102 7112 7158 7168
rect 6734 4528 6790 4584
rect 7572 13626 7628 13628
rect 7652 13626 7708 13628
rect 7732 13626 7788 13628
rect 7812 13626 7868 13628
rect 7572 13574 7618 13626
rect 7618 13574 7628 13626
rect 7652 13574 7682 13626
rect 7682 13574 7694 13626
rect 7694 13574 7708 13626
rect 7732 13574 7746 13626
rect 7746 13574 7758 13626
rect 7758 13574 7788 13626
rect 7812 13574 7822 13626
rect 7822 13574 7868 13626
rect 7572 13572 7628 13574
rect 7652 13572 7708 13574
rect 7732 13572 7788 13574
rect 7812 13572 7868 13574
rect 7470 13232 7526 13288
rect 8114 14728 8170 14784
rect 8942 14456 8998 14512
rect 8206 14048 8262 14104
rect 7930 13096 7986 13152
rect 7572 12538 7628 12540
rect 7652 12538 7708 12540
rect 7732 12538 7788 12540
rect 7812 12538 7868 12540
rect 7572 12486 7618 12538
rect 7618 12486 7628 12538
rect 7652 12486 7682 12538
rect 7682 12486 7694 12538
rect 7694 12486 7708 12538
rect 7732 12486 7746 12538
rect 7746 12486 7758 12538
rect 7758 12486 7788 12538
rect 7812 12486 7822 12538
rect 7822 12486 7868 12538
rect 7572 12484 7628 12486
rect 7652 12484 7708 12486
rect 7732 12484 7788 12486
rect 7812 12484 7868 12486
rect 7572 11450 7628 11452
rect 7652 11450 7708 11452
rect 7732 11450 7788 11452
rect 7812 11450 7868 11452
rect 7572 11398 7618 11450
rect 7618 11398 7628 11450
rect 7652 11398 7682 11450
rect 7682 11398 7694 11450
rect 7694 11398 7708 11450
rect 7732 11398 7746 11450
rect 7746 11398 7758 11450
rect 7758 11398 7788 11450
rect 7812 11398 7822 11450
rect 7822 11398 7868 11450
rect 7572 11396 7628 11398
rect 7652 11396 7708 11398
rect 7732 11396 7788 11398
rect 7812 11396 7868 11398
rect 7194 6024 7250 6080
rect 8206 13640 8262 13696
rect 8572 14170 8628 14172
rect 8652 14170 8708 14172
rect 8732 14170 8788 14172
rect 8812 14170 8868 14172
rect 8572 14118 8618 14170
rect 8618 14118 8628 14170
rect 8652 14118 8682 14170
rect 8682 14118 8694 14170
rect 8694 14118 8708 14170
rect 8732 14118 8746 14170
rect 8746 14118 8758 14170
rect 8758 14118 8788 14170
rect 8812 14118 8822 14170
rect 8822 14118 8868 14170
rect 8572 14116 8628 14118
rect 8652 14116 8708 14118
rect 8732 14116 8788 14118
rect 8812 14116 8868 14118
rect 8942 13812 8944 13832
rect 8944 13812 8996 13832
rect 8996 13812 8998 13832
rect 8942 13776 8998 13812
rect 8206 12824 8262 12880
rect 8206 12552 8262 12608
rect 8572 13082 8628 13084
rect 8652 13082 8708 13084
rect 8732 13082 8788 13084
rect 8812 13082 8868 13084
rect 8572 13030 8618 13082
rect 8618 13030 8628 13082
rect 8652 13030 8682 13082
rect 8682 13030 8694 13082
rect 8694 13030 8708 13082
rect 8732 13030 8746 13082
rect 8746 13030 8758 13082
rect 8758 13030 8788 13082
rect 8812 13030 8822 13082
rect 8822 13030 8868 13082
rect 8572 13028 8628 13030
rect 8652 13028 8708 13030
rect 8732 13028 8788 13030
rect 8812 13028 8868 13030
rect 8758 12280 8814 12336
rect 8572 11994 8628 11996
rect 8652 11994 8708 11996
rect 8732 11994 8788 11996
rect 8812 11994 8868 11996
rect 8572 11942 8618 11994
rect 8618 11942 8628 11994
rect 8652 11942 8682 11994
rect 8682 11942 8694 11994
rect 8694 11942 8708 11994
rect 8732 11942 8746 11994
rect 8746 11942 8758 11994
rect 8758 11942 8788 11994
rect 8812 11942 8822 11994
rect 8822 11942 8868 11994
rect 8572 11940 8628 11942
rect 8652 11940 8708 11942
rect 8732 11940 8788 11942
rect 8812 11940 8868 11942
rect 11058 15408 11114 15464
rect 9126 15308 9128 15328
rect 9128 15308 9180 15328
rect 9180 15308 9182 15328
rect 9126 15272 9182 15308
rect 9126 14320 9182 14376
rect 9126 14068 9182 14104
rect 9126 14048 9128 14068
rect 9128 14048 9180 14068
rect 9180 14048 9182 14068
rect 9310 14220 9312 14240
rect 9312 14220 9364 14240
rect 9364 14220 9366 14240
rect 9310 14184 9366 14220
rect 9218 12960 9274 13016
rect 12346 14456 12402 14512
rect 10782 14048 10838 14104
rect 11058 14048 11114 14104
rect 9678 13504 9734 13560
rect 9034 11736 9090 11792
rect 8758 11464 8814 11520
rect 8390 10784 8446 10840
rect 8390 10668 8446 10704
rect 8390 10648 8392 10668
rect 8392 10648 8444 10668
rect 8444 10648 8446 10668
rect 7572 10362 7628 10364
rect 7652 10362 7708 10364
rect 7732 10362 7788 10364
rect 7812 10362 7868 10364
rect 7572 10310 7618 10362
rect 7618 10310 7628 10362
rect 7652 10310 7682 10362
rect 7682 10310 7694 10362
rect 7694 10310 7708 10362
rect 7732 10310 7746 10362
rect 7746 10310 7758 10362
rect 7758 10310 7788 10362
rect 7812 10310 7822 10362
rect 7822 10310 7868 10362
rect 7572 10308 7628 10310
rect 7652 10308 7708 10310
rect 7732 10308 7788 10310
rect 7812 10308 7868 10310
rect 8022 9968 8078 10024
rect 7572 9274 7628 9276
rect 7652 9274 7708 9276
rect 7732 9274 7788 9276
rect 7812 9274 7868 9276
rect 7572 9222 7618 9274
rect 7618 9222 7628 9274
rect 7652 9222 7682 9274
rect 7682 9222 7694 9274
rect 7694 9222 7708 9274
rect 7732 9222 7746 9274
rect 7746 9222 7758 9274
rect 7758 9222 7788 9274
rect 7812 9222 7822 9274
rect 7822 9222 7868 9274
rect 7572 9220 7628 9222
rect 7652 9220 7708 9222
rect 7732 9220 7788 9222
rect 7812 9220 7868 9222
rect 7572 8186 7628 8188
rect 7652 8186 7708 8188
rect 7732 8186 7788 8188
rect 7812 8186 7868 8188
rect 7572 8134 7618 8186
rect 7618 8134 7628 8186
rect 7652 8134 7682 8186
rect 7682 8134 7694 8186
rect 7694 8134 7708 8186
rect 7732 8134 7746 8186
rect 7746 8134 7758 8186
rect 7758 8134 7788 8186
rect 7812 8134 7822 8186
rect 7822 8134 7868 8186
rect 7572 8132 7628 8134
rect 7652 8132 7708 8134
rect 7732 8132 7788 8134
rect 7812 8132 7868 8134
rect 7470 7928 7526 7984
rect 7572 7098 7628 7100
rect 7652 7098 7708 7100
rect 7732 7098 7788 7100
rect 7812 7098 7868 7100
rect 7572 7046 7618 7098
rect 7618 7046 7628 7098
rect 7652 7046 7682 7098
rect 7682 7046 7694 7098
rect 7694 7046 7708 7098
rect 7732 7046 7746 7098
rect 7746 7046 7758 7098
rect 7758 7046 7788 7098
rect 7812 7046 7822 7098
rect 7822 7046 7868 7098
rect 7572 7044 7628 7046
rect 7652 7044 7708 7046
rect 7732 7044 7788 7046
rect 7812 7044 7868 7046
rect 7286 4800 7342 4856
rect 7286 4392 7342 4448
rect 7010 3576 7066 3632
rect 6550 2932 6552 2952
rect 6552 2932 6604 2952
rect 6604 2932 6606 2952
rect 6550 2896 6606 2932
rect 5998 1672 6054 1728
rect 6182 1400 6238 1456
rect 6642 2488 6698 2544
rect 6734 2080 6790 2136
rect 7194 3440 7250 3496
rect 7572 6010 7628 6012
rect 7652 6010 7708 6012
rect 7732 6010 7788 6012
rect 7812 6010 7868 6012
rect 7572 5958 7618 6010
rect 7618 5958 7628 6010
rect 7652 5958 7682 6010
rect 7682 5958 7694 6010
rect 7694 5958 7708 6010
rect 7732 5958 7746 6010
rect 7746 5958 7758 6010
rect 7758 5958 7788 6010
rect 7812 5958 7822 6010
rect 7822 5958 7868 6010
rect 7572 5956 7628 5958
rect 7652 5956 7708 5958
rect 7732 5956 7788 5958
rect 7812 5956 7868 5958
rect 7746 5752 7802 5808
rect 7572 4922 7628 4924
rect 7652 4922 7708 4924
rect 7732 4922 7788 4924
rect 7812 4922 7868 4924
rect 7572 4870 7618 4922
rect 7618 4870 7628 4922
rect 7652 4870 7682 4922
rect 7682 4870 7694 4922
rect 7694 4870 7708 4922
rect 7732 4870 7746 4922
rect 7746 4870 7758 4922
rect 7758 4870 7788 4922
rect 7812 4870 7822 4922
rect 7822 4870 7868 4922
rect 7572 4868 7628 4870
rect 7652 4868 7708 4870
rect 7732 4868 7788 4870
rect 7812 4868 7868 4870
rect 7572 3834 7628 3836
rect 7652 3834 7708 3836
rect 7732 3834 7788 3836
rect 7812 3834 7868 3836
rect 7572 3782 7618 3834
rect 7618 3782 7628 3834
rect 7652 3782 7682 3834
rect 7682 3782 7694 3834
rect 7694 3782 7708 3834
rect 7732 3782 7746 3834
rect 7746 3782 7758 3834
rect 7758 3782 7788 3834
rect 7812 3782 7822 3834
rect 7822 3782 7868 3834
rect 7572 3780 7628 3782
rect 7652 3780 7708 3782
rect 7732 3780 7788 3782
rect 7812 3780 7868 3782
rect 7930 3304 7986 3360
rect 8298 9696 8354 9752
rect 8206 9152 8262 9208
rect 8114 5888 8170 5944
rect 8572 10906 8628 10908
rect 8652 10906 8708 10908
rect 8732 10906 8788 10908
rect 8812 10906 8868 10908
rect 8572 10854 8618 10906
rect 8618 10854 8628 10906
rect 8652 10854 8682 10906
rect 8682 10854 8694 10906
rect 8694 10854 8708 10906
rect 8732 10854 8746 10906
rect 8746 10854 8758 10906
rect 8758 10854 8788 10906
rect 8812 10854 8822 10906
rect 8822 10854 8868 10906
rect 8572 10852 8628 10854
rect 8652 10852 8708 10854
rect 8732 10852 8788 10854
rect 8812 10852 8868 10854
rect 8572 9818 8628 9820
rect 8652 9818 8708 9820
rect 8732 9818 8788 9820
rect 8812 9818 8868 9820
rect 8572 9766 8618 9818
rect 8618 9766 8628 9818
rect 8652 9766 8682 9818
rect 8682 9766 8694 9818
rect 8694 9766 8708 9818
rect 8732 9766 8746 9818
rect 8746 9766 8758 9818
rect 8758 9766 8788 9818
rect 8812 9766 8822 9818
rect 8822 9766 8868 9818
rect 8572 9764 8628 9766
rect 8652 9764 8708 9766
rect 8732 9764 8788 9766
rect 8812 9764 8868 9766
rect 8482 9560 8538 9616
rect 9310 11328 9366 11384
rect 9126 10648 9182 10704
rect 9494 10376 9550 10432
rect 10322 13096 10378 13152
rect 9862 11600 9918 11656
rect 10322 11056 10378 11112
rect 9862 10920 9918 10976
rect 10506 10648 10562 10704
rect 8572 8730 8628 8732
rect 8652 8730 8708 8732
rect 8732 8730 8788 8732
rect 8812 8730 8868 8732
rect 8572 8678 8618 8730
rect 8618 8678 8628 8730
rect 8652 8678 8682 8730
rect 8682 8678 8694 8730
rect 8694 8678 8708 8730
rect 8732 8678 8746 8730
rect 8746 8678 8758 8730
rect 8758 8678 8788 8730
rect 8812 8678 8822 8730
rect 8822 8678 8868 8730
rect 8572 8676 8628 8678
rect 8652 8676 8708 8678
rect 8732 8676 8788 8678
rect 8812 8676 8868 8678
rect 8390 7248 8446 7304
rect 8572 7642 8628 7644
rect 8652 7642 8708 7644
rect 8732 7642 8788 7644
rect 8812 7642 8868 7644
rect 8572 7590 8618 7642
rect 8618 7590 8628 7642
rect 8652 7590 8682 7642
rect 8682 7590 8694 7642
rect 8694 7590 8708 7642
rect 8732 7590 8746 7642
rect 8746 7590 8758 7642
rect 8758 7590 8788 7642
rect 8812 7590 8822 7642
rect 8822 7590 8868 7642
rect 8572 7588 8628 7590
rect 8652 7588 8708 7590
rect 8732 7588 8788 7590
rect 8812 7588 8868 7590
rect 9126 8336 9182 8392
rect 8482 6704 8538 6760
rect 8206 5364 8262 5400
rect 8206 5344 8208 5364
rect 8208 5344 8260 5364
rect 8260 5344 8262 5364
rect 8206 4392 8262 4448
rect 8572 6554 8628 6556
rect 8652 6554 8708 6556
rect 8732 6554 8788 6556
rect 8812 6554 8868 6556
rect 8572 6502 8618 6554
rect 8618 6502 8628 6554
rect 8652 6502 8682 6554
rect 8682 6502 8694 6554
rect 8694 6502 8708 6554
rect 8732 6502 8746 6554
rect 8746 6502 8758 6554
rect 8758 6502 8788 6554
rect 8812 6502 8822 6554
rect 8822 6502 8868 6554
rect 8572 6500 8628 6502
rect 8652 6500 8708 6502
rect 8732 6500 8788 6502
rect 8812 6500 8868 6502
rect 8850 6296 8906 6352
rect 8572 5466 8628 5468
rect 8652 5466 8708 5468
rect 8732 5466 8788 5468
rect 8812 5466 8868 5468
rect 8572 5414 8618 5466
rect 8618 5414 8628 5466
rect 8652 5414 8682 5466
rect 8682 5414 8694 5466
rect 8694 5414 8708 5466
rect 8732 5414 8746 5466
rect 8746 5414 8758 5466
rect 8758 5414 8788 5466
rect 8812 5414 8822 5466
rect 8822 5414 8868 5466
rect 8572 5412 8628 5414
rect 8652 5412 8708 5414
rect 8732 5412 8788 5414
rect 8812 5412 8868 5414
rect 8572 4378 8628 4380
rect 8652 4378 8708 4380
rect 8732 4378 8788 4380
rect 8812 4378 8868 4380
rect 8572 4326 8618 4378
rect 8618 4326 8628 4378
rect 8652 4326 8682 4378
rect 8682 4326 8694 4378
rect 8694 4326 8708 4378
rect 8732 4326 8746 4378
rect 8746 4326 8758 4378
rect 8758 4326 8788 4378
rect 8812 4326 8822 4378
rect 8822 4326 8868 4378
rect 8572 4324 8628 4326
rect 8652 4324 8708 4326
rect 8732 4324 8788 4326
rect 8812 4324 8868 4326
rect 8206 3712 8262 3768
rect 7572 2746 7628 2748
rect 7652 2746 7708 2748
rect 7732 2746 7788 2748
rect 7812 2746 7868 2748
rect 7572 2694 7618 2746
rect 7618 2694 7628 2746
rect 7652 2694 7682 2746
rect 7682 2694 7694 2746
rect 7694 2694 7708 2746
rect 7732 2694 7746 2746
rect 7746 2694 7758 2746
rect 7758 2694 7788 2746
rect 7812 2694 7822 2746
rect 7822 2694 7868 2746
rect 7572 2692 7628 2694
rect 7652 2692 7708 2694
rect 7732 2692 7788 2694
rect 7812 2692 7868 2694
rect 9310 7404 9366 7440
rect 9310 7384 9312 7404
rect 9312 7384 9364 7404
rect 9364 7384 9366 7404
rect 8572 3290 8628 3292
rect 8652 3290 8708 3292
rect 8732 3290 8788 3292
rect 8812 3290 8868 3292
rect 8572 3238 8618 3290
rect 8618 3238 8628 3290
rect 8652 3238 8682 3290
rect 8682 3238 8694 3290
rect 8694 3238 8708 3290
rect 8732 3238 8746 3290
rect 8746 3238 8758 3290
rect 8758 3238 8788 3290
rect 8812 3238 8822 3290
rect 8822 3238 8868 3290
rect 8572 3236 8628 3238
rect 8652 3236 8708 3238
rect 8732 3236 8788 3238
rect 8812 3236 8868 3238
rect 8298 3168 8354 3224
rect 9126 4664 9182 4720
rect 9218 3884 9220 3904
rect 9220 3884 9272 3904
rect 9272 3884 9274 3904
rect 9218 3848 9274 3884
rect 9218 3440 9274 3496
rect 9126 3168 9182 3224
rect 9034 2896 9090 2952
rect 9218 2916 9274 2952
rect 9218 2896 9220 2916
rect 9220 2896 9272 2916
rect 9272 2896 9274 2916
rect 8758 2760 8814 2816
rect 9218 2624 9274 2680
rect 8758 2352 8814 2408
rect 8942 2352 8998 2408
rect 7470 1828 7526 1864
rect 7470 1808 7472 1828
rect 7472 1808 7524 1828
rect 7524 1808 7526 1828
rect 7572 1658 7628 1660
rect 7652 1658 7708 1660
rect 7732 1658 7788 1660
rect 7812 1658 7868 1660
rect 7572 1606 7618 1658
rect 7618 1606 7628 1658
rect 7652 1606 7682 1658
rect 7682 1606 7694 1658
rect 7694 1606 7708 1658
rect 7732 1606 7746 1658
rect 7746 1606 7758 1658
rect 7758 1606 7788 1658
rect 7812 1606 7822 1658
rect 7822 1606 7868 1658
rect 7572 1604 7628 1606
rect 7652 1604 7708 1606
rect 7732 1604 7788 1606
rect 7812 1604 7868 1606
rect 3606 1300 3608 1320
rect 3608 1300 3660 1320
rect 3660 1300 3662 1320
rect 3606 1264 3662 1300
rect 4066 1284 4122 1320
rect 7378 1300 7380 1320
rect 7380 1300 7432 1320
rect 7432 1300 7434 1320
rect 4066 1264 4068 1284
rect 4068 1264 4120 1284
rect 4120 1264 4122 1284
rect 2870 1128 2926 1184
rect 3572 1114 3628 1116
rect 3652 1114 3708 1116
rect 3732 1114 3788 1116
rect 3812 1114 3868 1116
rect 3572 1062 3618 1114
rect 3618 1062 3628 1114
rect 3652 1062 3682 1114
rect 3682 1062 3694 1114
rect 3694 1062 3708 1114
rect 3732 1062 3746 1114
rect 3746 1062 3758 1114
rect 3758 1062 3788 1114
rect 3812 1062 3822 1114
rect 3822 1062 3868 1114
rect 3572 1060 3628 1062
rect 3652 1060 3708 1062
rect 3732 1060 3788 1062
rect 3812 1060 3868 1062
rect 1030 856 1086 912
rect 5998 992 6054 1048
rect 4894 856 4950 912
rect 4342 720 4398 776
rect 4158 584 4214 640
rect 7378 1264 7434 1300
rect 8206 1284 8262 1320
rect 8206 1264 8208 1284
rect 8208 1264 8260 1284
rect 8260 1264 8262 1284
rect 8390 2216 8446 2272
rect 8572 2202 8628 2204
rect 8652 2202 8708 2204
rect 8732 2202 8788 2204
rect 8812 2202 8868 2204
rect 8572 2150 8618 2202
rect 8618 2150 8628 2202
rect 8652 2150 8682 2202
rect 8682 2150 8694 2202
rect 8694 2150 8708 2202
rect 8732 2150 8746 2202
rect 8746 2150 8758 2202
rect 8758 2150 8788 2202
rect 8812 2150 8822 2202
rect 8822 2150 8868 2202
rect 8572 2148 8628 2150
rect 8652 2148 8708 2150
rect 8732 2148 8788 2150
rect 8812 2148 8868 2150
rect 9034 2216 9090 2272
rect 8390 1672 8446 1728
rect 8572 1114 8628 1116
rect 8652 1114 8708 1116
rect 8732 1114 8788 1116
rect 8812 1114 8868 1116
rect 8572 1062 8618 1114
rect 8618 1062 8628 1114
rect 8652 1062 8682 1114
rect 8682 1062 8694 1114
rect 8694 1062 8708 1114
rect 8732 1062 8746 1114
rect 8746 1062 8758 1114
rect 8758 1062 8788 1114
rect 8812 1062 8822 1114
rect 8822 1062 8868 1114
rect 8572 1060 8628 1062
rect 8652 1060 8708 1062
rect 8732 1060 8788 1062
rect 8812 1060 8868 1062
rect 8114 584 8170 640
rect 8298 584 8354 640
rect 6734 312 6790 368
rect 9402 5480 9458 5536
rect 9770 9016 9826 9072
rect 9770 4936 9826 4992
rect 9770 3576 9826 3632
rect 9954 5364 10010 5400
rect 9954 5344 9956 5364
rect 9956 5344 10008 5364
rect 10008 5344 10010 5364
rect 9954 3596 10010 3632
rect 9954 3576 9956 3596
rect 9956 3576 10008 3596
rect 10008 3576 10010 3596
rect 11058 13776 11114 13832
rect 10966 8200 11022 8256
rect 10966 5888 11022 5944
rect 12806 14204 12862 14240
rect 12806 14184 12808 14204
rect 12808 14184 12860 14204
rect 12860 14184 12862 14204
rect 12438 13912 12494 13968
rect 12346 13232 12402 13288
rect 12346 12824 12402 12880
rect 11150 6432 11206 6488
rect 11058 5616 11114 5672
rect 11150 5208 11206 5264
rect 11058 5072 11114 5128
rect 11058 3304 11114 3360
rect 10874 2896 10930 2952
rect 9310 2080 9366 2136
rect 9586 2080 9642 2136
rect 11702 7792 11758 7848
rect 11518 6568 11574 6624
rect 11334 5752 11390 5808
rect 11886 6976 11942 7032
rect 11794 6024 11850 6080
rect 11702 5480 11758 5536
rect 11518 3440 11574 3496
rect 12806 12008 12862 12064
rect 12714 11328 12770 11384
rect 12530 10920 12586 10976
rect 12622 9968 12678 10024
rect 12530 6432 12586 6488
rect 12346 6160 12402 6216
rect 11886 4528 11942 4584
rect 12070 4528 12126 4584
rect 11702 3304 11758 3360
rect 11242 1808 11298 1864
rect 12254 3168 12310 3224
rect 12714 4800 12770 4856
rect 12622 3712 12678 3768
rect 12898 11464 12954 11520
rect 12806 3576 12862 3632
rect 13450 15952 13506 16008
rect 13450 12824 13506 12880
rect 13450 12708 13506 12744
rect 13450 12688 13452 12708
rect 13452 12688 13504 12708
rect 13504 12688 13506 12708
rect 13634 15952 13690 16008
rect 13634 15292 13690 15328
rect 13634 15272 13636 15292
rect 13636 15272 13688 15292
rect 13688 15272 13690 15292
rect 13634 14884 13690 14920
rect 13634 14864 13636 14884
rect 13636 14864 13688 14884
rect 13688 14864 13690 14884
rect 13634 14748 13690 14784
rect 13634 14728 13636 14748
rect 13636 14728 13688 14748
rect 13688 14728 13690 14748
rect 13634 14612 13690 14648
rect 13634 14592 13636 14612
rect 13636 14592 13688 14612
rect 13688 14592 13690 14612
rect 17912 15544 17968 15600
rect 13818 14764 13820 14784
rect 13820 14764 13872 14784
rect 13872 14764 13874 14784
rect 13818 14728 13874 14764
rect 13726 14320 13782 14376
rect 13634 14184 13690 14240
rect 13542 11484 13598 11520
rect 13542 11464 13544 11484
rect 13544 11464 13596 11484
rect 13596 11464 13598 11484
rect 13726 13640 13782 13696
rect 13818 13524 13874 13560
rect 13818 13504 13820 13524
rect 13820 13504 13872 13524
rect 13872 13504 13874 13524
rect 13726 13368 13782 13424
rect 13818 12980 13874 13016
rect 13818 12960 13820 12980
rect 13820 12960 13872 12980
rect 13872 12960 13874 12980
rect 13818 12572 13874 12608
rect 13818 12552 13820 12572
rect 13820 12552 13872 12572
rect 13872 12552 13874 12572
rect 13818 12180 13820 12200
rect 13820 12180 13872 12200
rect 13872 12180 13874 12200
rect 13818 12144 13874 12180
rect 13818 11908 13820 11928
rect 13820 11908 13872 11928
rect 13872 11908 13874 11928
rect 13818 11872 13874 11908
rect 13818 11192 13874 11248
rect 13634 10648 13690 10704
rect 13542 10512 13598 10568
rect 13174 9460 13176 9480
rect 13176 9460 13228 9480
rect 13228 9460 13230 9480
rect 13174 9424 13230 9460
rect 13450 9152 13506 9208
rect 13266 6024 13322 6080
rect 13818 10376 13874 10432
rect 13818 10276 13820 10296
rect 13820 10276 13872 10296
rect 13872 10276 13874 10296
rect 13818 10240 13874 10276
rect 13726 9696 13782 9752
rect 13818 9288 13874 9344
rect 13818 9052 13820 9072
rect 13820 9052 13872 9072
rect 13872 9052 13874 9072
rect 13818 9016 13874 9052
rect 13818 7420 13820 7440
rect 13820 7420 13872 7440
rect 13872 7420 13874 7440
rect 13818 7384 13874 7420
rect 13818 6840 13874 6896
rect 13818 5788 13820 5808
rect 13820 5788 13872 5808
rect 13872 5788 13874 5808
rect 13818 5752 13874 5788
rect 13634 5244 13636 5264
rect 13636 5244 13688 5264
rect 13688 5244 13690 5264
rect 13634 5208 13690 5244
rect 13818 5344 13874 5400
rect 13726 5072 13782 5128
rect 13450 4936 13506 4992
rect 13726 4800 13782 4856
rect 13726 4120 13782 4176
rect 13818 3712 13874 3768
rect 12990 3304 13046 3360
rect 12346 2760 12402 2816
rect 12070 2216 12126 2272
rect 13818 1944 13874 2000
rect 11702 1672 11758 1728
rect 9126 448 9182 504
rect 13910 312 13966 368
rect 17912 15156 17968 15192
rect 17912 15136 17914 15156
rect 17914 15136 17966 15156
rect 17966 15136 17968 15156
rect 16854 2352 16910 2408
rect 17314 4120 17370 4176
rect 17912 13540 17914 13560
rect 17914 13540 17966 13560
rect 17966 13540 17968 13560
rect 17912 13504 17968 13540
rect 17912 6180 17968 6216
rect 17912 6160 17914 6180
rect 17914 6160 17966 6180
rect 17966 6160 17968 6180
rect 18050 3848 18106 3904
rect 18050 2488 18106 2544
rect 16946 1536 17002 1592
rect 15106 1400 15162 1456
rect 14278 856 14334 912
rect 19062 16632 19118 16688
rect 18326 3712 18382 3768
rect 18418 2080 18474 2136
rect 17774 720 17830 776
rect 18510 1264 18566 1320
rect 17866 584 17922 640
rect 18786 4256 18842 4312
rect 18970 3984 19026 4040
rect 19062 3032 19118 3088
rect 18602 448 18658 504
rect 8114 176 8170 232
rect 14094 176 14150 232
<< metal3 >>
rect 2405 16962 2471 16965
rect 18413 16962 18479 16965
rect 2405 16960 18479 16962
rect 2405 16904 2410 16960
rect 2466 16904 18418 16960
rect 18474 16904 18479 16960
rect 2405 16902 18479 16904
rect 2405 16899 2471 16902
rect 18413 16899 18479 16902
rect 3141 16826 3207 16829
rect 13629 16826 13695 16829
rect 3141 16824 13695 16826
rect 3141 16768 3146 16824
rect 3202 16768 13634 16824
rect 13690 16768 13695 16824
rect 3141 16766 13695 16768
rect 3141 16763 3207 16766
rect 13629 16763 13695 16766
rect 4705 16690 4771 16693
rect 13721 16690 13787 16693
rect 15101 16690 15167 16693
rect 4705 16688 13787 16690
rect 4705 16632 4710 16688
rect 4766 16632 13726 16688
rect 13782 16632 13787 16688
rect 4705 16630 13787 16632
rect 4705 16627 4771 16630
rect 13721 16627 13787 16630
rect 13862 16688 15167 16690
rect 13862 16632 15106 16688
rect 15162 16632 15167 16688
rect 13862 16630 15167 16632
rect 6177 16282 6243 16285
rect 13862 16282 13922 16630
rect 15101 16627 15167 16630
rect 15285 16690 15351 16693
rect 18229 16690 18295 16693
rect 19057 16690 19123 16693
rect 15285 16688 18295 16690
rect 15285 16632 15290 16688
rect 15346 16632 18234 16688
rect 18290 16632 18295 16688
rect 15285 16630 18295 16632
rect 15285 16627 15351 16630
rect 18229 16627 18295 16630
rect 19014 16688 19123 16690
rect 19014 16632 19062 16688
rect 19118 16632 19123 16688
rect 19014 16627 19123 16632
rect 19014 16448 19074 16627
rect 14000 16328 34000 16448
rect 6177 16280 13922 16282
rect 6177 16224 6182 16280
rect 6238 16224 13922 16280
rect 6177 16222 13922 16224
rect 6177 16219 6243 16222
rect 4061 16146 4127 16149
rect 13077 16146 13143 16149
rect 4061 16144 13143 16146
rect 4061 16088 4066 16144
rect 4122 16088 13082 16144
rect 13138 16088 13143 16144
rect 4061 16086 13143 16088
rect 4061 16083 4127 16086
rect 13077 16083 13143 16086
rect 5717 16010 5783 16013
rect 13445 16010 13511 16013
rect 5717 16008 13511 16010
rect 5717 15952 5722 16008
rect 5778 15952 13450 16008
rect 13506 15952 13511 16008
rect 5717 15950 13511 15952
rect 5717 15947 5783 15950
rect 13445 15947 13511 15950
rect 13629 16010 13695 16013
rect 14000 16010 34000 16040
rect 13629 16008 34000 16010
rect 13629 15952 13634 16008
rect 13690 15952 34000 16008
rect 13629 15950 34000 15952
rect 13629 15947 13695 15950
rect 14000 15920 34000 15950
rect 2562 15808 2878 15809
rect 2562 15744 2568 15808
rect 2632 15744 2648 15808
rect 2712 15744 2728 15808
rect 2792 15744 2808 15808
rect 2872 15744 2878 15808
rect 2562 15743 2878 15744
rect 7562 15808 7878 15809
rect 7562 15744 7568 15808
rect 7632 15744 7648 15808
rect 7712 15744 7728 15808
rect 7792 15744 7808 15808
rect 7872 15744 7878 15808
rect 7562 15743 7878 15744
rect 14000 15600 34000 15632
rect 14000 15544 17912 15600
rect 17968 15544 34000 15600
rect 14000 15512 34000 15544
rect 1761 15466 1827 15469
rect 5257 15466 5323 15469
rect 1761 15464 5323 15466
rect 1761 15408 1766 15464
rect 1822 15408 5262 15464
rect 5318 15408 5323 15464
rect 1761 15406 5323 15408
rect 1761 15403 1827 15406
rect 5257 15403 5323 15406
rect 8109 15466 8175 15469
rect 11053 15466 11119 15469
rect 8109 15464 11119 15466
rect 8109 15408 8114 15464
rect 8170 15408 11058 15464
rect 11114 15408 11119 15464
rect 8109 15406 11119 15408
rect 8109 15403 8175 15406
rect 11053 15403 11119 15406
rect 381 15330 447 15333
rect 2773 15330 2839 15333
rect 381 15328 2839 15330
rect 381 15272 386 15328
rect 442 15272 2778 15328
rect 2834 15272 2839 15328
rect 381 15270 2839 15272
rect 381 15267 447 15270
rect 2773 15267 2839 15270
rect 9121 15330 9187 15333
rect 13629 15330 13695 15333
rect 9121 15328 13695 15330
rect 9121 15272 9126 15328
rect 9182 15272 13634 15328
rect 13690 15272 13695 15328
rect 9121 15270 13695 15272
rect 9121 15267 9187 15270
rect 13629 15267 13695 15270
rect 3562 15264 3878 15265
rect 3562 15200 3568 15264
rect 3632 15200 3648 15264
rect 3712 15200 3728 15264
rect 3792 15200 3808 15264
rect 3872 15200 3878 15264
rect 3562 15199 3878 15200
rect 8562 15264 8878 15265
rect 8562 15200 8568 15264
rect 8632 15200 8648 15264
rect 8712 15200 8728 15264
rect 8792 15200 8808 15264
rect 8872 15200 8878 15264
rect 8562 15199 8878 15200
rect 6545 15194 6611 15197
rect 8385 15194 8451 15197
rect 6545 15192 8451 15194
rect 6545 15136 6550 15192
rect 6606 15136 8390 15192
rect 8446 15136 8451 15192
rect 6545 15134 8451 15136
rect 6545 15131 6611 15134
rect 8385 15131 8451 15134
rect 14000 15192 34000 15224
rect 14000 15136 17912 15192
rect 17968 15136 34000 15192
rect 14000 15104 34000 15136
rect 4061 15058 4127 15061
rect 5349 15058 5415 15061
rect 4061 15056 5415 15058
rect 4061 15000 4066 15056
rect 4122 15000 5354 15056
rect 5410 15000 5415 15056
rect 4061 14998 5415 15000
rect 4061 14995 4127 14998
rect 5349 14995 5415 14998
rect 473 14922 539 14925
rect 2773 14922 2839 14925
rect 473 14920 2839 14922
rect 473 14864 478 14920
rect 534 14864 2778 14920
rect 2834 14864 2839 14920
rect 473 14862 2839 14864
rect 473 14859 539 14862
rect 2773 14859 2839 14862
rect 5441 14922 5507 14925
rect 13629 14922 13695 14925
rect 5441 14920 13695 14922
rect 5441 14864 5446 14920
rect 5502 14864 13634 14920
rect 13690 14864 13695 14920
rect 5441 14862 13695 14864
rect 5441 14859 5507 14862
rect 13629 14859 13695 14862
rect 8109 14786 8175 14789
rect 13629 14786 13695 14789
rect 8109 14784 13695 14786
rect 8109 14728 8114 14784
rect 8170 14728 13634 14784
rect 13690 14728 13695 14784
rect 8109 14726 13695 14728
rect 8109 14723 8175 14726
rect 13629 14723 13695 14726
rect 13813 14786 13879 14789
rect 14000 14786 34000 14816
rect 13813 14784 34000 14786
rect 13813 14728 13818 14784
rect 13874 14728 34000 14784
rect 13813 14726 34000 14728
rect 13813 14723 13879 14726
rect 2562 14720 2878 14721
rect 2562 14656 2568 14720
rect 2632 14656 2648 14720
rect 2712 14656 2728 14720
rect 2792 14656 2808 14720
rect 2872 14656 2878 14720
rect 2562 14655 2878 14656
rect 7562 14720 7878 14721
rect 7562 14656 7568 14720
rect 7632 14656 7648 14720
rect 7712 14656 7728 14720
rect 7792 14656 7808 14720
rect 7872 14656 7878 14720
rect 14000 14696 34000 14726
rect 7562 14655 7878 14656
rect 13629 14650 13695 14653
rect 8342 14648 13695 14650
rect 8342 14592 13634 14648
rect 13690 14592 13695 14648
rect 8342 14590 13695 14592
rect 197 14514 263 14517
rect 4429 14514 4495 14517
rect 197 14512 4495 14514
rect 197 14456 202 14512
rect 258 14456 4434 14512
rect 4490 14456 4495 14512
rect 197 14454 4495 14456
rect 197 14451 263 14454
rect 4429 14451 4495 14454
rect 3969 14378 4035 14381
rect 6913 14378 6979 14381
rect 3969 14376 6979 14378
rect 3969 14320 3974 14376
rect 4030 14320 6918 14376
rect 6974 14320 6979 14376
rect 3969 14318 6979 14320
rect 3969 14315 4035 14318
rect 6913 14315 6979 14318
rect 4061 14242 4127 14245
rect 8342 14242 8402 14590
rect 13629 14587 13695 14590
rect 8937 14514 9003 14517
rect 12341 14514 12407 14517
rect 8937 14512 12407 14514
rect 8937 14456 8942 14512
rect 8998 14456 12346 14512
rect 12402 14456 12407 14512
rect 8937 14454 12407 14456
rect 8937 14451 9003 14454
rect 12341 14451 12407 14454
rect 9121 14378 9187 14381
rect 13721 14378 13787 14381
rect 14000 14378 34000 14408
rect 9121 14376 13002 14378
rect 9121 14320 9126 14376
rect 9182 14320 13002 14376
rect 9121 14318 13002 14320
rect 9121 14315 9187 14318
rect 4061 14240 8402 14242
rect 4061 14184 4066 14240
rect 4122 14184 8402 14240
rect 4061 14182 8402 14184
rect 9305 14242 9371 14245
rect 12801 14242 12867 14245
rect 9305 14240 12867 14242
rect 9305 14184 9310 14240
rect 9366 14184 12806 14240
rect 12862 14184 12867 14240
rect 9305 14182 12867 14184
rect 12942 14242 13002 14318
rect 13721 14376 34000 14378
rect 13721 14320 13726 14376
rect 13782 14320 34000 14376
rect 13721 14318 34000 14320
rect 13721 14315 13787 14318
rect 14000 14288 34000 14318
rect 13629 14242 13695 14245
rect 12942 14240 13695 14242
rect 12942 14184 13634 14240
rect 13690 14184 13695 14240
rect 12942 14182 13695 14184
rect 4061 14179 4127 14182
rect 9305 14179 9371 14182
rect 12801 14179 12867 14182
rect 13629 14179 13695 14182
rect 3562 14176 3878 14177
rect 3562 14112 3568 14176
rect 3632 14112 3648 14176
rect 3712 14112 3728 14176
rect 3792 14112 3808 14176
rect 3872 14112 3878 14176
rect 3562 14111 3878 14112
rect 8562 14176 8878 14177
rect 8562 14112 8568 14176
rect 8632 14112 8648 14176
rect 8712 14112 8728 14176
rect 8792 14112 8808 14176
rect 8872 14112 8878 14176
rect 8562 14111 8878 14112
rect 4061 14106 4127 14109
rect 8201 14106 8267 14109
rect 4061 14104 8267 14106
rect 4061 14048 4066 14104
rect 4122 14048 8206 14104
rect 8262 14048 8267 14104
rect 4061 14046 8267 14048
rect 4061 14043 4127 14046
rect 8201 14043 8267 14046
rect 9121 14106 9187 14109
rect 10777 14106 10843 14109
rect 9121 14104 10843 14106
rect 9121 14048 9126 14104
rect 9182 14048 10782 14104
rect 10838 14048 10843 14104
rect 9121 14046 10843 14048
rect 9121 14043 9187 14046
rect 10777 14043 10843 14046
rect 11053 14106 11119 14109
rect 11053 14104 13186 14106
rect 11053 14048 11058 14104
rect 11114 14048 13186 14104
rect 11053 14046 13186 14048
rect 11053 14043 11119 14046
rect 2497 13970 2563 13973
rect 3141 13970 3207 13973
rect 2497 13968 3207 13970
rect 2497 13912 2502 13968
rect 2558 13912 3146 13968
rect 3202 13912 3207 13968
rect 2497 13910 3207 13912
rect 2497 13907 2563 13910
rect 3141 13907 3207 13910
rect 4889 13970 4955 13973
rect 12433 13970 12499 13973
rect 4889 13968 12499 13970
rect 4889 13912 4894 13968
rect 4950 13912 12438 13968
rect 12494 13912 12499 13968
rect 4889 13910 12499 13912
rect 13126 13970 13186 14046
rect 14000 13970 34000 14000
rect 13126 13910 34000 13970
rect 4889 13907 4955 13910
rect 12433 13907 12499 13910
rect 14000 13880 34000 13910
rect 1209 13834 1275 13837
rect 2773 13834 2839 13837
rect 1209 13832 2839 13834
rect 1209 13776 1214 13832
rect 1270 13776 2778 13832
rect 2834 13776 2839 13832
rect 1209 13774 2839 13776
rect 1209 13771 1275 13774
rect 2773 13771 2839 13774
rect 6637 13834 6703 13837
rect 7230 13834 7236 13836
rect 6637 13832 7236 13834
rect 6637 13776 6642 13832
rect 6698 13776 7236 13832
rect 6637 13774 7236 13776
rect 6637 13771 6703 13774
rect 7230 13772 7236 13774
rect 7300 13772 7306 13836
rect 8937 13834 9003 13837
rect 11053 13834 11119 13837
rect 7422 13774 8034 13834
rect 2562 13632 2878 13633
rect 2562 13568 2568 13632
rect 2632 13568 2648 13632
rect 2712 13568 2728 13632
rect 2792 13568 2808 13632
rect 2872 13568 2878 13632
rect 2562 13567 2878 13568
rect 7422 13562 7482 13774
rect 7562 13632 7878 13633
rect 7562 13568 7568 13632
rect 7632 13568 7648 13632
rect 7712 13568 7728 13632
rect 7792 13568 7808 13632
rect 7872 13568 7878 13632
rect 7562 13567 7878 13568
rect 6870 13502 7482 13562
rect 7974 13562 8034 13774
rect 8937 13832 11119 13834
rect 8937 13776 8942 13832
rect 8998 13776 11058 13832
rect 11114 13776 11119 13832
rect 8937 13774 11119 13776
rect 8937 13771 9003 13774
rect 11053 13771 11119 13774
rect 8201 13698 8267 13701
rect 13721 13698 13787 13701
rect 8201 13696 13787 13698
rect 8201 13640 8206 13696
rect 8262 13640 13726 13696
rect 13782 13640 13787 13696
rect 8201 13638 13787 13640
rect 8201 13635 8267 13638
rect 13721 13635 13787 13638
rect 9673 13562 9739 13565
rect 13813 13562 13879 13565
rect 7974 13560 9739 13562
rect 7974 13504 9678 13560
rect 9734 13504 9739 13560
rect 7974 13502 9739 13504
rect 3417 13426 3483 13429
rect 6870 13426 6930 13502
rect 9673 13499 9739 13502
rect 12390 13560 13879 13562
rect 12390 13504 13818 13560
rect 13874 13504 13879 13560
rect 12390 13502 13879 13504
rect 3417 13424 6930 13426
rect 3417 13368 3422 13424
rect 3478 13368 6930 13424
rect 3417 13366 6930 13368
rect 7005 13426 7071 13429
rect 12390 13426 12450 13502
rect 13813 13499 13879 13502
rect 14000 13560 34000 13592
rect 14000 13504 17912 13560
rect 17968 13504 34000 13560
rect 14000 13472 34000 13504
rect 13721 13426 13787 13429
rect 7005 13424 12450 13426
rect 7005 13368 7010 13424
rect 7066 13368 12450 13424
rect 7005 13366 12450 13368
rect 13126 13424 13787 13426
rect 13126 13368 13726 13424
rect 13782 13368 13787 13424
rect 13126 13366 13787 13368
rect 3417 13363 3483 13366
rect 7005 13363 7071 13366
rect 2221 13290 2287 13293
rect 7465 13290 7531 13293
rect 2221 13288 7531 13290
rect 2221 13232 2226 13288
rect 2282 13232 7470 13288
rect 7526 13232 7531 13288
rect 2221 13230 7531 13232
rect 2221 13227 2287 13230
rect 7465 13227 7531 13230
rect 12341 13290 12407 13293
rect 13126 13290 13186 13366
rect 13721 13363 13787 13366
rect 12341 13288 13186 13290
rect 12341 13232 12346 13288
rect 12402 13232 13186 13288
rect 12341 13230 13186 13232
rect 12341 13227 12407 13230
rect 4061 13154 4127 13157
rect 7925 13154 7991 13157
rect 4061 13152 7991 13154
rect 4061 13096 4066 13152
rect 4122 13096 7930 13152
rect 7986 13096 7991 13152
rect 4061 13094 7991 13096
rect 4061 13091 4127 13094
rect 7925 13091 7991 13094
rect 10317 13154 10383 13157
rect 14000 13154 34000 13184
rect 10317 13152 34000 13154
rect 10317 13096 10322 13152
rect 10378 13096 34000 13152
rect 10317 13094 34000 13096
rect 10317 13091 10383 13094
rect 3562 13088 3878 13089
rect 3562 13024 3568 13088
rect 3632 13024 3648 13088
rect 3712 13024 3728 13088
rect 3792 13024 3808 13088
rect 3872 13024 3878 13088
rect 3562 13023 3878 13024
rect 8562 13088 8878 13089
rect 8562 13024 8568 13088
rect 8632 13024 8648 13088
rect 8712 13024 8728 13088
rect 8792 13024 8808 13088
rect 8872 13024 8878 13088
rect 14000 13064 34000 13094
rect 8562 13023 8878 13024
rect 4429 13018 4495 13021
rect 9213 13018 9279 13021
rect 13813 13018 13879 13021
rect 4429 13016 8402 13018
rect 4429 12960 4434 13016
rect 4490 12960 8402 13016
rect 4429 12958 8402 12960
rect 4429 12955 4495 12958
rect 6637 12882 6703 12885
rect 8201 12882 8267 12885
rect 6637 12880 8267 12882
rect 6637 12824 6642 12880
rect 6698 12824 8206 12880
rect 8262 12824 8267 12880
rect 6637 12822 8267 12824
rect 8342 12882 8402 12958
rect 9213 13016 13879 13018
rect 9213 12960 9218 13016
rect 9274 12960 13818 13016
rect 13874 12960 13879 13016
rect 9213 12958 13879 12960
rect 9213 12955 9279 12958
rect 13813 12955 13879 12958
rect 12341 12882 12407 12885
rect 8342 12880 12407 12882
rect 8342 12824 12346 12880
rect 12402 12824 12407 12880
rect 8342 12822 12407 12824
rect 6637 12819 6703 12822
rect 8201 12819 8267 12822
rect 12341 12819 12407 12822
rect 13445 12882 13511 12885
rect 13445 12880 13922 12882
rect 13445 12824 13450 12880
rect 13506 12824 13922 12880
rect 13445 12822 13922 12824
rect 13445 12819 13511 12822
rect 2589 12746 2655 12749
rect 13445 12746 13511 12749
rect 2589 12744 13511 12746
rect 2589 12688 2594 12744
rect 2650 12688 13450 12744
rect 13506 12688 13511 12744
rect 2589 12686 13511 12688
rect 13862 12746 13922 12822
rect 14000 12746 34000 12776
rect 13862 12686 34000 12746
rect 2589 12683 2655 12686
rect 13445 12683 13511 12686
rect 14000 12656 34000 12686
rect 8201 12610 8267 12613
rect 13813 12610 13879 12613
rect 8201 12608 13879 12610
rect 8201 12552 8206 12608
rect 8262 12552 13818 12608
rect 13874 12552 13879 12608
rect 8201 12550 13879 12552
rect 8201 12547 8267 12550
rect 13813 12547 13879 12550
rect 2562 12544 2878 12545
rect 2562 12480 2568 12544
rect 2632 12480 2648 12544
rect 2712 12480 2728 12544
rect 2792 12480 2808 12544
rect 2872 12480 2878 12544
rect 2562 12479 2878 12480
rect 7562 12544 7878 12545
rect 7562 12480 7568 12544
rect 7632 12480 7648 12544
rect 7712 12480 7728 12544
rect 7792 12480 7808 12544
rect 7872 12480 7878 12544
rect 7562 12479 7878 12480
rect 1577 12474 1643 12477
rect 1350 12472 1643 12474
rect 1350 12416 1582 12472
rect 1638 12416 1643 12472
rect 1350 12414 1643 12416
rect 1350 12340 1410 12414
rect 1577 12411 1643 12414
rect 1342 12276 1348 12340
rect 1412 12276 1418 12340
rect 6085 12338 6151 12341
rect 8753 12338 8819 12341
rect 14000 12338 34000 12368
rect 6085 12336 8819 12338
rect 6085 12280 6090 12336
rect 6146 12280 8758 12336
rect 8814 12280 8819 12336
rect 6085 12278 8819 12280
rect 6085 12275 6151 12278
rect 8753 12275 8819 12278
rect 13862 12278 34000 12338
rect 13862 12205 13922 12278
rect 14000 12248 34000 12278
rect 565 12202 631 12205
rect 3509 12202 3575 12205
rect 565 12200 3575 12202
rect 565 12144 570 12200
rect 626 12144 3514 12200
rect 3570 12144 3575 12200
rect 565 12142 3575 12144
rect 565 12139 631 12142
rect 3509 12139 3575 12142
rect 5993 12202 6059 12205
rect 5993 12200 12450 12202
rect 5993 12144 5998 12200
rect 6054 12144 12450 12200
rect 5993 12142 12450 12144
rect 5993 12139 6059 12142
rect 1301 12068 1367 12069
rect 1301 12064 1348 12068
rect 1412 12066 1418 12068
rect 12390 12066 12450 12142
rect 13813 12200 13922 12205
rect 13813 12144 13818 12200
rect 13874 12144 13922 12200
rect 13813 12142 13922 12144
rect 13813 12139 13879 12142
rect 12801 12066 12867 12069
rect 1301 12008 1306 12064
rect 1301 12004 1348 12008
rect 1412 12006 1458 12066
rect 12390 12064 12867 12066
rect 12390 12008 12806 12064
rect 12862 12008 12867 12064
rect 12390 12006 12867 12008
rect 1412 12004 1418 12006
rect 1301 12003 1367 12004
rect 12801 12003 12867 12006
rect 3562 12000 3878 12001
rect 3562 11936 3568 12000
rect 3632 11936 3648 12000
rect 3712 11936 3728 12000
rect 3792 11936 3808 12000
rect 3872 11936 3878 12000
rect 3562 11935 3878 11936
rect 8562 12000 8878 12001
rect 8562 11936 8568 12000
rect 8632 11936 8648 12000
rect 8712 11936 8728 12000
rect 8792 11936 8808 12000
rect 8872 11936 8878 12000
rect 8562 11935 8878 11936
rect 4337 11930 4403 11933
rect 13813 11930 13879 11933
rect 14000 11930 34000 11960
rect 4337 11928 8402 11930
rect 4337 11872 4342 11928
rect 4398 11872 8402 11928
rect 4337 11870 8402 11872
rect 4337 11867 4403 11870
rect 2129 11794 2195 11797
rect 5533 11794 5599 11797
rect 2129 11792 5599 11794
rect 2129 11736 2134 11792
rect 2190 11736 5538 11792
rect 5594 11736 5599 11792
rect 2129 11734 5599 11736
rect 8342 11794 8402 11870
rect 13813 11928 34000 11930
rect 13813 11872 13818 11928
rect 13874 11872 34000 11928
rect 13813 11870 34000 11872
rect 13813 11867 13879 11870
rect 14000 11840 34000 11870
rect 9029 11794 9095 11797
rect 8342 11792 9095 11794
rect 8342 11736 9034 11792
rect 9090 11736 9095 11792
rect 8342 11734 9095 11736
rect 2129 11731 2195 11734
rect 5533 11731 5599 11734
rect 9029 11731 9095 11734
rect 1393 11658 1459 11661
rect 4153 11658 4219 11661
rect 1393 11656 4219 11658
rect 1393 11600 1398 11656
rect 1454 11600 4158 11656
rect 4214 11600 4219 11656
rect 1393 11598 4219 11600
rect 1393 11595 1459 11598
rect 4153 11595 4219 11598
rect 6269 11658 6335 11661
rect 9857 11658 9923 11661
rect 6269 11656 9923 11658
rect 6269 11600 6274 11656
rect 6330 11600 9862 11656
rect 9918 11600 9923 11656
rect 6269 11598 9923 11600
rect 6269 11595 6335 11598
rect 9857 11595 9923 11598
rect 3601 11522 3667 11525
rect 4889 11522 4955 11525
rect 6361 11522 6427 11525
rect 3601 11520 6427 11522
rect 3601 11464 3606 11520
rect 3662 11464 4894 11520
rect 4950 11464 6366 11520
rect 6422 11464 6427 11520
rect 3601 11462 6427 11464
rect 3601 11459 3667 11462
rect 4889 11459 4955 11462
rect 6361 11459 6427 11462
rect 8753 11522 8819 11525
rect 12893 11522 12959 11525
rect 8753 11520 12959 11522
rect 8753 11464 8758 11520
rect 8814 11464 12898 11520
rect 12954 11464 12959 11520
rect 8753 11462 12959 11464
rect 8753 11459 8819 11462
rect 12893 11459 12959 11462
rect 13537 11522 13603 11525
rect 14000 11522 34000 11552
rect 13537 11520 34000 11522
rect 13537 11464 13542 11520
rect 13598 11464 34000 11520
rect 13537 11462 34000 11464
rect 13537 11459 13603 11462
rect 2562 11456 2878 11457
rect 2562 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2878 11456
rect 2562 11391 2878 11392
rect 7562 11456 7878 11457
rect 7562 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7878 11456
rect 14000 11432 34000 11462
rect 7562 11391 7878 11392
rect 6085 11386 6151 11389
rect 5214 11384 6151 11386
rect 5214 11328 6090 11384
rect 6146 11328 6151 11384
rect 5214 11326 6151 11328
rect 2681 11250 2747 11253
rect 5214 11250 5274 11326
rect 6085 11323 6151 11326
rect 9305 11386 9371 11389
rect 12709 11386 12775 11389
rect 9305 11384 12775 11386
rect 9305 11328 9310 11384
rect 9366 11328 12714 11384
rect 12770 11328 12775 11384
rect 9305 11326 12775 11328
rect 9305 11323 9371 11326
rect 12709 11323 12775 11326
rect 2681 11248 5274 11250
rect 2681 11192 2686 11248
rect 2742 11192 5274 11248
rect 2681 11190 5274 11192
rect 5441 11250 5507 11253
rect 7097 11250 7163 11253
rect 5441 11248 7163 11250
rect 5441 11192 5446 11248
rect 5502 11192 7102 11248
rect 7158 11192 7163 11248
rect 5441 11190 7163 11192
rect 2681 11187 2747 11190
rect 5441 11187 5507 11190
rect 7097 11187 7163 11190
rect 13813 11250 13879 11253
rect 13813 11248 13922 11250
rect 13813 11192 13818 11248
rect 13874 11192 13922 11248
rect 13813 11187 13922 11192
rect 933 11114 999 11117
rect 3233 11114 3299 11117
rect 933 11112 3299 11114
rect 933 11056 938 11112
rect 994 11056 3238 11112
rect 3294 11056 3299 11112
rect 933 11054 3299 11056
rect 933 11051 999 11054
rect 3233 11051 3299 11054
rect 4061 11114 4127 11117
rect 4981 11114 5047 11117
rect 6453 11114 6519 11117
rect 4061 11112 4170 11114
rect 4061 11056 4066 11112
rect 4122 11056 4170 11112
rect 4061 11051 4170 11056
rect 4981 11112 6519 11114
rect 4981 11056 4986 11112
rect 5042 11056 6458 11112
rect 6514 11056 6519 11112
rect 4981 11054 6519 11056
rect 4981 11051 5047 11054
rect 6453 11051 6519 11054
rect 7189 11114 7255 11117
rect 10317 11114 10383 11117
rect 7189 11112 10383 11114
rect 7189 11056 7194 11112
rect 7250 11056 10322 11112
rect 10378 11056 10383 11112
rect 7189 11054 10383 11056
rect 13862 11114 13922 11187
rect 14000 11114 34000 11144
rect 13862 11054 34000 11114
rect 7189 11051 7255 11054
rect 10317 11051 10383 11054
rect 4110 10978 4170 11051
rect 14000 11024 34000 11054
rect 7005 10978 7071 10981
rect 4110 10976 7071 10978
rect 4110 10920 7010 10976
rect 7066 10920 7071 10976
rect 4110 10918 7071 10920
rect 7005 10915 7071 10918
rect 9857 10978 9923 10981
rect 12525 10978 12591 10981
rect 9857 10976 12591 10978
rect 9857 10920 9862 10976
rect 9918 10920 12530 10976
rect 12586 10920 12591 10976
rect 9857 10918 12591 10920
rect 9857 10915 9923 10918
rect 12525 10915 12591 10918
rect 3562 10912 3878 10913
rect 3562 10848 3568 10912
rect 3632 10848 3648 10912
rect 3712 10848 3728 10912
rect 3792 10848 3808 10912
rect 3872 10848 3878 10912
rect 3562 10847 3878 10848
rect 8562 10912 8878 10913
rect 8562 10848 8568 10912
rect 8632 10848 8648 10912
rect 8712 10848 8728 10912
rect 8792 10848 8808 10912
rect 8872 10848 8878 10912
rect 8562 10847 8878 10848
rect 4797 10842 4863 10845
rect 8385 10842 8451 10845
rect 4797 10840 8451 10842
rect 4797 10784 4802 10840
rect 4858 10784 8390 10840
rect 8446 10784 8451 10840
rect 4797 10782 8451 10784
rect 4797 10779 4863 10782
rect 8385 10779 8451 10782
rect 6913 10706 6979 10709
rect 8385 10706 8451 10709
rect 6913 10704 8451 10706
rect 6913 10648 6918 10704
rect 6974 10648 8390 10704
rect 8446 10648 8451 10704
rect 6913 10646 8451 10648
rect 6913 10643 6979 10646
rect 8385 10643 8451 10646
rect 9121 10706 9187 10709
rect 10501 10706 10567 10709
rect 9121 10704 10567 10706
rect 9121 10648 9126 10704
rect 9182 10648 10506 10704
rect 10562 10648 10567 10704
rect 9121 10646 10567 10648
rect 9121 10643 9187 10646
rect 10501 10643 10567 10646
rect 13629 10706 13695 10709
rect 14000 10706 34000 10736
rect 13629 10704 34000 10706
rect 13629 10648 13634 10704
rect 13690 10648 34000 10704
rect 13629 10646 34000 10648
rect 13629 10643 13695 10646
rect 14000 10616 34000 10646
rect 2497 10570 2563 10573
rect 13537 10570 13603 10573
rect 2497 10568 13603 10570
rect 2497 10512 2502 10568
rect 2558 10512 13542 10568
rect 13598 10512 13603 10568
rect 2497 10510 13603 10512
rect 2497 10507 2563 10510
rect 13537 10507 13603 10510
rect 9489 10434 9555 10437
rect 13813 10434 13879 10437
rect 9489 10432 13879 10434
rect 9489 10376 9494 10432
rect 9550 10376 13818 10432
rect 13874 10376 13879 10432
rect 9489 10374 13879 10376
rect 9489 10371 9555 10374
rect 13813 10371 13879 10374
rect 2562 10368 2878 10369
rect 2562 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2878 10368
rect 2562 10303 2878 10304
rect 7562 10368 7878 10369
rect 7562 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7878 10368
rect 7562 10303 7878 10304
rect 13813 10298 13879 10301
rect 14000 10298 34000 10328
rect 13813 10296 34000 10298
rect 13813 10240 13818 10296
rect 13874 10240 34000 10296
rect 13813 10238 34000 10240
rect 13813 10235 13879 10238
rect 14000 10208 34000 10238
rect 2957 10162 3023 10165
rect 7097 10162 7163 10165
rect 2957 10160 7163 10162
rect 2957 10104 2962 10160
rect 3018 10104 7102 10160
rect 7158 10104 7163 10160
rect 2957 10102 7163 10104
rect 2957 10099 3023 10102
rect 7097 10099 7163 10102
rect 3325 10026 3391 10029
rect 4337 10026 4403 10029
rect 3325 10024 4403 10026
rect 3325 9968 3330 10024
rect 3386 9968 4342 10024
rect 4398 9968 4403 10024
rect 3325 9966 4403 9968
rect 3325 9963 3391 9966
rect 4337 9963 4403 9966
rect 8017 10026 8083 10029
rect 12617 10026 12683 10029
rect 8017 10024 12683 10026
rect 8017 9968 8022 10024
rect 8078 9968 12622 10024
rect 12678 9968 12683 10024
rect 8017 9966 12683 9968
rect 8017 9963 8083 9966
rect 12617 9963 12683 9966
rect 14000 9890 34000 9920
rect 13862 9830 34000 9890
rect 3562 9824 3878 9825
rect 3562 9760 3568 9824
rect 3632 9760 3648 9824
rect 3712 9760 3728 9824
rect 3792 9760 3808 9824
rect 3872 9760 3878 9824
rect 3562 9759 3878 9760
rect 8562 9824 8878 9825
rect 8562 9760 8568 9824
rect 8632 9760 8648 9824
rect 8712 9760 8728 9824
rect 8792 9760 8808 9824
rect 8872 9760 8878 9824
rect 8562 9759 8878 9760
rect 749 9754 815 9757
rect 3233 9754 3299 9757
rect 749 9752 3299 9754
rect 749 9696 754 9752
rect 810 9696 3238 9752
rect 3294 9696 3299 9752
rect 749 9694 3299 9696
rect 749 9691 815 9694
rect 3233 9691 3299 9694
rect 4521 9754 4587 9757
rect 5625 9754 5691 9757
rect 4521 9752 5691 9754
rect 4521 9696 4526 9752
rect 4582 9696 5630 9752
rect 5686 9696 5691 9752
rect 4521 9694 5691 9696
rect 4521 9691 4587 9694
rect 5625 9691 5691 9694
rect 5993 9754 6059 9757
rect 8293 9754 8359 9757
rect 5993 9752 8359 9754
rect 5993 9696 5998 9752
rect 6054 9696 8298 9752
rect 8354 9696 8359 9752
rect 5993 9694 8359 9696
rect 5993 9691 6059 9694
rect 8293 9691 8359 9694
rect 13721 9754 13787 9757
rect 13862 9754 13922 9830
rect 14000 9800 34000 9830
rect 13721 9752 13922 9754
rect 13721 9696 13726 9752
rect 13782 9696 13922 9752
rect 13721 9694 13922 9696
rect 13721 9691 13787 9694
rect 5809 9618 5875 9621
rect 8477 9618 8543 9621
rect 5809 9616 8543 9618
rect 5809 9560 5814 9616
rect 5870 9560 8482 9616
rect 8538 9560 8543 9616
rect 5809 9558 8543 9560
rect 5809 9555 5875 9558
rect 8477 9555 8543 9558
rect 2681 9482 2747 9485
rect 13169 9482 13235 9485
rect 14000 9482 34000 9512
rect 2681 9480 13235 9482
rect 2681 9424 2686 9480
rect 2742 9424 13174 9480
rect 13230 9424 13235 9480
rect 2681 9422 13235 9424
rect 2681 9419 2747 9422
rect 13169 9419 13235 9422
rect 13862 9422 34000 9482
rect 13862 9349 13922 9422
rect 14000 9392 34000 9422
rect 5993 9346 6059 9349
rect 7230 9346 7236 9348
rect 5993 9344 7236 9346
rect 5993 9288 5998 9344
rect 6054 9288 7236 9344
rect 5993 9286 7236 9288
rect 5993 9283 6059 9286
rect 7230 9284 7236 9286
rect 7300 9284 7306 9348
rect 13813 9344 13922 9349
rect 13813 9288 13818 9344
rect 13874 9288 13922 9344
rect 13813 9286 13922 9288
rect 2562 9280 2878 9281
rect 2562 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2878 9280
rect 2562 9215 2878 9216
rect 4061 9210 4127 9213
rect 5809 9210 5875 9213
rect 4061 9208 5875 9210
rect 4061 9152 4066 9208
rect 4122 9152 5814 9208
rect 5870 9152 5875 9208
rect 4061 9150 5875 9152
rect 4061 9147 4127 9150
rect 5809 9147 5875 9150
rect 1117 9074 1183 9077
rect 4981 9074 5047 9077
rect 1117 9072 5047 9074
rect 1117 9016 1122 9072
rect 1178 9016 4986 9072
rect 5042 9016 5047 9072
rect 1117 9014 5047 9016
rect 7238 9074 7298 9284
rect 13813 9283 13879 9286
rect 7562 9280 7878 9281
rect 7562 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7878 9280
rect 7562 9215 7878 9216
rect 8201 9210 8267 9213
rect 13445 9210 13511 9213
rect 8201 9208 13511 9210
rect 8201 9152 8206 9208
rect 8262 9152 13450 9208
rect 13506 9152 13511 9208
rect 8201 9150 13511 9152
rect 8201 9147 8267 9150
rect 13445 9147 13511 9150
rect 9765 9074 9831 9077
rect 7238 9072 9831 9074
rect 7238 9016 9770 9072
rect 9826 9016 9831 9072
rect 7238 9014 9831 9016
rect 1117 9011 1183 9014
rect 4981 9011 5047 9014
rect 9765 9011 9831 9014
rect 13813 9074 13879 9077
rect 14000 9074 34000 9104
rect 13813 9072 34000 9074
rect 13813 9016 13818 9072
rect 13874 9016 34000 9072
rect 13813 9014 34000 9016
rect 13813 9011 13879 9014
rect 14000 8984 34000 9014
rect 3233 8938 3299 8941
rect 8334 8938 8340 8940
rect 3233 8936 8340 8938
rect 3233 8880 3238 8936
rect 3294 8880 8340 8936
rect 3233 8878 8340 8880
rect 3233 8875 3299 8878
rect 8334 8876 8340 8878
rect 8404 8876 8410 8940
rect 3562 8736 3878 8737
rect 3562 8672 3568 8736
rect 3632 8672 3648 8736
rect 3712 8672 3728 8736
rect 3792 8672 3808 8736
rect 3872 8672 3878 8736
rect 3562 8671 3878 8672
rect 8562 8736 8878 8737
rect 8562 8672 8568 8736
rect 8632 8672 8648 8736
rect 8712 8672 8728 8736
rect 8792 8672 8808 8736
rect 8872 8672 8878 8736
rect 8562 8671 8878 8672
rect 14000 8666 34000 8696
rect 12390 8606 34000 8666
rect 5625 8530 5691 8533
rect 12390 8530 12450 8606
rect 14000 8576 34000 8606
rect 5625 8528 12450 8530
rect 5625 8472 5630 8528
rect 5686 8472 12450 8528
rect 5625 8470 12450 8472
rect 5625 8467 5691 8470
rect 1117 8394 1183 8397
rect 2773 8394 2839 8397
rect 1117 8392 2839 8394
rect 1117 8336 1122 8392
rect 1178 8336 2778 8392
rect 2834 8336 2839 8392
rect 1117 8334 2839 8336
rect 1117 8331 1183 8334
rect 2773 8331 2839 8334
rect 5349 8394 5415 8397
rect 9121 8394 9187 8397
rect 5349 8392 9187 8394
rect 5349 8336 5354 8392
rect 5410 8336 9126 8392
rect 9182 8336 9187 8392
rect 5349 8334 9187 8336
rect 5349 8331 5415 8334
rect 9121 8331 9187 8334
rect 10961 8258 11027 8261
rect 14000 8258 34000 8288
rect 10961 8256 34000 8258
rect 10961 8200 10966 8256
rect 11022 8200 34000 8256
rect 10961 8198 34000 8200
rect 10961 8195 11027 8198
rect 2562 8192 2878 8193
rect 2562 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2878 8192
rect 2562 8127 2878 8128
rect 7562 8192 7878 8193
rect 7562 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7878 8192
rect 14000 8168 34000 8198
rect 7562 8127 7878 8128
rect 2405 7986 2471 7989
rect 3049 7986 3115 7989
rect 2405 7984 3115 7986
rect 2405 7928 2410 7984
rect 2466 7928 3054 7984
rect 3110 7928 3115 7984
rect 2405 7926 3115 7928
rect 2405 7923 2471 7926
rect 3049 7923 3115 7926
rect 3877 7986 3943 7989
rect 7465 7986 7531 7989
rect 3877 7984 7531 7986
rect 3877 7928 3882 7984
rect 3938 7928 7470 7984
rect 7526 7928 7531 7984
rect 3877 7926 7531 7928
rect 3877 7923 3943 7926
rect 7465 7923 7531 7926
rect 1025 7850 1091 7853
rect 3509 7850 3575 7853
rect 1025 7848 3575 7850
rect 1025 7792 1030 7848
rect 1086 7792 3514 7848
rect 3570 7792 3575 7848
rect 1025 7790 3575 7792
rect 1025 7787 1091 7790
rect 3509 7787 3575 7790
rect 11697 7850 11763 7853
rect 14000 7850 34000 7880
rect 11697 7848 34000 7850
rect 11697 7792 11702 7848
rect 11758 7792 34000 7848
rect 11697 7790 34000 7792
rect 11697 7787 11763 7790
rect 14000 7760 34000 7790
rect 3562 7648 3878 7649
rect 3562 7584 3568 7648
rect 3632 7584 3648 7648
rect 3712 7584 3728 7648
rect 3792 7584 3808 7648
rect 3872 7584 3878 7648
rect 3562 7583 3878 7584
rect 8562 7648 8878 7649
rect 8562 7584 8568 7648
rect 8632 7584 8648 7648
rect 8712 7584 8728 7648
rect 8792 7584 8808 7648
rect 8872 7584 8878 7648
rect 8562 7583 8878 7584
rect 2221 7442 2287 7445
rect 9305 7442 9371 7445
rect 2221 7440 9371 7442
rect 2221 7384 2226 7440
rect 2282 7384 9310 7440
rect 9366 7384 9371 7440
rect 2221 7382 9371 7384
rect 2221 7379 2287 7382
rect 9305 7379 9371 7382
rect 13813 7442 13879 7445
rect 14000 7442 34000 7472
rect 13813 7440 34000 7442
rect 13813 7384 13818 7440
rect 13874 7384 34000 7440
rect 13813 7382 34000 7384
rect 13813 7379 13879 7382
rect 14000 7352 34000 7382
rect 3233 7306 3299 7309
rect 8385 7306 8451 7309
rect 3233 7304 8451 7306
rect 3233 7248 3238 7304
rect 3294 7248 8390 7304
rect 8446 7248 8451 7304
rect 3233 7246 8451 7248
rect 3233 7243 3299 7246
rect 8385 7243 8451 7246
rect 5349 7170 5415 7173
rect 7097 7170 7163 7173
rect 5349 7168 7163 7170
rect 5349 7112 5354 7168
rect 5410 7112 7102 7168
rect 7158 7112 7163 7168
rect 5349 7110 7163 7112
rect 5349 7107 5415 7110
rect 7097 7107 7163 7110
rect 2562 7104 2878 7105
rect 2562 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2878 7104
rect 2562 7039 2878 7040
rect 7562 7104 7878 7105
rect 7562 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7878 7104
rect 7562 7039 7878 7040
rect 4061 7034 4127 7037
rect 6361 7034 6427 7037
rect 4061 7032 6427 7034
rect 4061 6976 4066 7032
rect 4122 6976 6366 7032
rect 6422 6976 6427 7032
rect 4061 6974 6427 6976
rect 4061 6971 4127 6974
rect 6361 6971 6427 6974
rect 11881 7034 11947 7037
rect 14000 7034 34000 7064
rect 11881 7032 34000 7034
rect 11881 6976 11886 7032
rect 11942 6976 34000 7032
rect 11881 6974 34000 6976
rect 11881 6971 11947 6974
rect 14000 6944 34000 6974
rect 1577 6898 1643 6901
rect 3049 6898 3115 6901
rect 13813 6898 13879 6901
rect 1577 6896 2790 6898
rect 1577 6840 1582 6896
rect 1638 6840 2790 6896
rect 1577 6838 2790 6840
rect 1577 6835 1643 6838
rect 2730 6762 2790 6838
rect 3049 6896 13879 6898
rect 3049 6840 3054 6896
rect 3110 6840 13818 6896
rect 13874 6840 13879 6896
rect 3049 6838 13879 6840
rect 3049 6835 3115 6838
rect 13813 6835 13879 6838
rect 4521 6762 4587 6765
rect 2730 6760 4587 6762
rect 2730 6704 4526 6760
rect 4582 6704 4587 6760
rect 2730 6702 4587 6704
rect 4521 6699 4587 6702
rect 6637 6762 6703 6765
rect 8477 6762 8543 6765
rect 6637 6760 8543 6762
rect 6637 6704 6642 6760
rect 6698 6704 8482 6760
rect 8538 6704 8543 6760
rect 6637 6702 8543 6704
rect 6637 6699 6703 6702
rect 8477 6699 8543 6702
rect 11513 6626 11579 6629
rect 14000 6626 34000 6656
rect 11513 6624 34000 6626
rect 11513 6568 11518 6624
rect 11574 6568 34000 6624
rect 11513 6566 34000 6568
rect 11513 6563 11579 6566
rect 3562 6560 3878 6561
rect 3562 6496 3568 6560
rect 3632 6496 3648 6560
rect 3712 6496 3728 6560
rect 3792 6496 3808 6560
rect 3872 6496 3878 6560
rect 3562 6495 3878 6496
rect 8562 6560 8878 6561
rect 8562 6496 8568 6560
rect 8632 6496 8648 6560
rect 8712 6496 8728 6560
rect 8792 6496 8808 6560
rect 8872 6496 8878 6560
rect 14000 6536 34000 6566
rect 8562 6495 8878 6496
rect 6269 6490 6335 6493
rect 11145 6490 11211 6493
rect 12525 6490 12591 6493
rect 6269 6488 8402 6490
rect 6269 6432 6274 6488
rect 6330 6432 8402 6488
rect 6269 6430 8402 6432
rect 6269 6427 6335 6430
rect 3509 6354 3575 6357
rect 6545 6354 6611 6357
rect 3509 6352 6611 6354
rect 3509 6296 3514 6352
rect 3570 6296 6550 6352
rect 6606 6296 6611 6352
rect 3509 6294 6611 6296
rect 8342 6354 8402 6430
rect 11145 6488 12591 6490
rect 11145 6432 11150 6488
rect 11206 6432 12530 6488
rect 12586 6432 12591 6488
rect 11145 6430 12591 6432
rect 11145 6427 11211 6430
rect 12525 6427 12591 6430
rect 8845 6354 8911 6357
rect 8342 6352 8911 6354
rect 8342 6296 8850 6352
rect 8906 6296 8911 6352
rect 8342 6294 8911 6296
rect 3509 6291 3575 6294
rect 6545 6291 6611 6294
rect 8845 6291 8911 6294
rect 5993 6218 6059 6221
rect 12341 6218 12407 6221
rect 5993 6216 12407 6218
rect 5993 6160 5998 6216
rect 6054 6160 12346 6216
rect 12402 6160 12407 6216
rect 5993 6158 12407 6160
rect 5993 6155 6059 6158
rect 12341 6155 12407 6158
rect 14000 6216 34000 6248
rect 14000 6160 17912 6216
rect 17968 6160 34000 6216
rect 14000 6128 34000 6160
rect 5441 6082 5507 6085
rect 7189 6082 7255 6085
rect 5441 6080 7255 6082
rect 5441 6024 5446 6080
rect 5502 6024 7194 6080
rect 7250 6024 7255 6080
rect 5441 6022 7255 6024
rect 5441 6019 5507 6022
rect 7189 6019 7255 6022
rect 11789 6082 11855 6085
rect 13261 6082 13327 6085
rect 11789 6080 13327 6082
rect 11789 6024 11794 6080
rect 11850 6024 13266 6080
rect 13322 6024 13327 6080
rect 11789 6022 13327 6024
rect 11789 6019 11855 6022
rect 13261 6019 13327 6022
rect 2562 6016 2878 6017
rect 2562 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2878 6016
rect 2562 5951 2878 5952
rect 7562 6016 7878 6017
rect 7562 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7878 6016
rect 7562 5951 7878 5952
rect 3049 5946 3115 5949
rect 4613 5946 4679 5949
rect 3049 5944 4679 5946
rect 3049 5888 3054 5944
rect 3110 5888 4618 5944
rect 4674 5888 4679 5944
rect 3049 5886 4679 5888
rect 3049 5883 3115 5886
rect 4613 5883 4679 5886
rect 8109 5946 8175 5949
rect 10961 5946 11027 5949
rect 8109 5944 11027 5946
rect 8109 5888 8114 5944
rect 8170 5888 10966 5944
rect 11022 5888 11027 5944
rect 8109 5886 11027 5888
rect 8109 5883 8175 5886
rect 10961 5883 11027 5886
rect 13816 5813 13922 5844
rect 4613 5810 4679 5813
rect 6177 5810 6243 5813
rect 4613 5808 6243 5810
rect 4613 5752 4618 5808
rect 4674 5752 6182 5808
rect 6238 5752 6243 5808
rect 4613 5750 6243 5752
rect 4613 5747 4679 5750
rect 6177 5747 6243 5750
rect 7741 5810 7807 5813
rect 11329 5810 11395 5813
rect 7741 5808 11395 5810
rect 7741 5752 7746 5808
rect 7802 5752 11334 5808
rect 11390 5752 11395 5808
rect 7741 5750 11395 5752
rect 7741 5747 7807 5750
rect 11329 5747 11395 5750
rect 13813 5810 13922 5813
rect 14000 5810 34000 5840
rect 13813 5808 34000 5810
rect 13813 5752 13818 5808
rect 13874 5752 34000 5808
rect 13813 5750 34000 5752
rect 13813 5747 13879 5750
rect 14000 5720 34000 5750
rect 2497 5674 2563 5677
rect 4797 5674 4863 5677
rect 2497 5672 4863 5674
rect 2497 5616 2502 5672
rect 2558 5616 4802 5672
rect 4858 5616 4863 5672
rect 2497 5614 4863 5616
rect 2497 5611 2563 5614
rect 4797 5611 4863 5614
rect 4981 5674 5047 5677
rect 11053 5674 11119 5677
rect 4981 5672 11119 5674
rect 4981 5616 4986 5672
rect 5042 5616 11058 5672
rect 11114 5616 11119 5672
rect 4981 5614 11119 5616
rect 4981 5611 5047 5614
rect 11053 5611 11119 5614
rect 9397 5538 9463 5541
rect 11697 5538 11763 5541
rect 9397 5536 11763 5538
rect 9397 5480 9402 5536
rect 9458 5480 11702 5536
rect 11758 5480 11763 5536
rect 9397 5478 11763 5480
rect 9397 5475 9463 5478
rect 11697 5475 11763 5478
rect 3562 5472 3878 5473
rect 3562 5408 3568 5472
rect 3632 5408 3648 5472
rect 3712 5408 3728 5472
rect 3792 5408 3808 5472
rect 3872 5408 3878 5472
rect 3562 5407 3878 5408
rect 8562 5472 8878 5473
rect 8562 5408 8568 5472
rect 8632 5408 8648 5472
rect 8712 5408 8728 5472
rect 8792 5408 8808 5472
rect 8872 5408 8878 5472
rect 8562 5407 8878 5408
rect 6361 5402 6427 5405
rect 8201 5402 8267 5405
rect 6361 5400 8267 5402
rect 6361 5344 6366 5400
rect 6422 5344 8206 5400
rect 8262 5344 8267 5400
rect 6361 5342 8267 5344
rect 6361 5339 6427 5342
rect 8201 5339 8267 5342
rect 9949 5402 10015 5405
rect 13813 5402 13879 5405
rect 14000 5402 34000 5432
rect 9949 5400 12450 5402
rect 9949 5344 9954 5400
rect 10010 5344 12450 5400
rect 9949 5342 12450 5344
rect 9949 5339 10015 5342
rect 1393 5266 1459 5269
rect 4521 5266 4587 5269
rect 1393 5264 4587 5266
rect 1393 5208 1398 5264
rect 1454 5208 4526 5264
rect 4582 5208 4587 5264
rect 1393 5206 4587 5208
rect 1393 5203 1459 5206
rect 4521 5203 4587 5206
rect 4705 5266 4771 5269
rect 11145 5266 11211 5269
rect 4705 5264 11211 5266
rect 4705 5208 4710 5264
rect 4766 5208 11150 5264
rect 11206 5208 11211 5264
rect 4705 5206 11211 5208
rect 12390 5266 12450 5342
rect 13813 5400 34000 5402
rect 13813 5344 13818 5400
rect 13874 5344 34000 5400
rect 13813 5342 34000 5344
rect 13813 5339 13879 5342
rect 14000 5312 34000 5342
rect 13629 5266 13695 5269
rect 12390 5264 13695 5266
rect 12390 5208 13634 5264
rect 13690 5208 13695 5264
rect 12390 5206 13695 5208
rect 4705 5203 4771 5206
rect 11145 5203 11211 5206
rect 13629 5203 13695 5206
rect 4153 5130 4219 5133
rect 11053 5130 11119 5133
rect 13721 5130 13787 5133
rect 4153 5128 8402 5130
rect 4153 5072 4158 5128
rect 4214 5072 8402 5128
rect 4153 5070 8402 5072
rect 4153 5067 4219 5070
rect 5441 4994 5507 4997
rect 5030 4992 5507 4994
rect 5030 4936 5446 4992
rect 5502 4936 5507 4992
rect 5030 4934 5507 4936
rect 2405 4858 2471 4861
rect 4889 4858 4955 4861
rect 2405 4856 4955 4858
rect 2405 4800 2410 4856
rect 2466 4800 4894 4856
rect 4950 4800 4955 4856
rect 2405 4798 4955 4800
rect 2405 4795 2471 4798
rect 4889 4795 4955 4798
rect 1301 4722 1367 4725
rect 3509 4722 3575 4725
rect 1301 4720 3575 4722
rect 1301 4664 1306 4720
rect 1362 4664 3514 4720
rect 3570 4664 3575 4720
rect 1301 4662 3575 4664
rect 1301 4659 1367 4662
rect 3509 4659 3575 4662
rect 4705 4722 4771 4725
rect 5030 4722 5090 4934
rect 5441 4931 5507 4934
rect 7562 4928 7878 4929
rect 7562 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7878 4928
rect 7562 4863 7878 4864
rect 5441 4858 5507 4861
rect 7281 4858 7347 4861
rect 5441 4856 7347 4858
rect 5441 4800 5446 4856
rect 5502 4800 7286 4856
rect 7342 4800 7347 4856
rect 5441 4798 7347 4800
rect 8342 4858 8402 5070
rect 11053 5128 13787 5130
rect 11053 5072 11058 5128
rect 11114 5072 13726 5128
rect 13782 5072 13787 5128
rect 11053 5070 13787 5072
rect 11053 5067 11119 5070
rect 13721 5067 13787 5070
rect 9765 4994 9831 4997
rect 13445 4994 13511 4997
rect 14000 4994 34000 5024
rect 9765 4992 13370 4994
rect 9765 4936 9770 4992
rect 9826 4936 13370 4992
rect 9765 4934 13370 4936
rect 9765 4931 9831 4934
rect 12709 4858 12775 4861
rect 8342 4856 12775 4858
rect 8342 4800 12714 4856
rect 12770 4800 12775 4856
rect 8342 4798 12775 4800
rect 13310 4858 13370 4934
rect 13445 4992 34000 4994
rect 13445 4936 13450 4992
rect 13506 4936 34000 4992
rect 13445 4934 34000 4936
rect 13445 4931 13511 4934
rect 14000 4904 34000 4934
rect 13721 4858 13787 4861
rect 13310 4856 13787 4858
rect 13310 4800 13726 4856
rect 13782 4800 13787 4856
rect 13310 4798 13787 4800
rect 5441 4795 5507 4798
rect 7281 4795 7347 4798
rect 12709 4795 12775 4798
rect 13721 4795 13787 4798
rect 4705 4720 5090 4722
rect 4705 4664 4710 4720
rect 4766 4664 5090 4720
rect 4705 4662 5090 4664
rect 6177 4722 6243 4725
rect 9121 4722 9187 4725
rect 6177 4720 9187 4722
rect 6177 4664 6182 4720
rect 6238 4664 9126 4720
rect 9182 4664 9187 4720
rect 6177 4662 9187 4664
rect 4705 4659 4771 4662
rect 6177 4659 6243 4662
rect 9121 4659 9187 4662
rect 6729 4586 6795 4589
rect 11881 4586 11947 4589
rect 6729 4584 11947 4586
rect 6729 4528 6734 4584
rect 6790 4528 11886 4584
rect 11942 4528 11947 4584
rect 6729 4526 11947 4528
rect 6729 4523 6795 4526
rect 11881 4523 11947 4526
rect 12065 4586 12131 4589
rect 14000 4586 34000 4616
rect 12065 4584 34000 4586
rect 12065 4528 12070 4584
rect 12126 4528 34000 4584
rect 12065 4526 34000 4528
rect 12065 4523 12131 4526
rect 14000 4496 34000 4526
rect 7281 4450 7347 4453
rect 8201 4450 8267 4453
rect 7281 4448 8267 4450
rect 7281 4392 7286 4448
rect 7342 4392 8206 4448
rect 8262 4392 8267 4448
rect 7281 4390 8267 4392
rect 7281 4387 7347 4390
rect 8201 4387 8267 4390
rect 3562 4384 3878 4385
rect 3562 4320 3568 4384
rect 3632 4320 3648 4384
rect 3712 4320 3728 4384
rect 3792 4320 3808 4384
rect 3872 4320 3878 4384
rect 3562 4319 3878 4320
rect 8562 4384 8878 4385
rect 8562 4320 8568 4384
rect 8632 4320 8648 4384
rect 8712 4320 8728 4384
rect 8792 4320 8808 4384
rect 8872 4320 8878 4384
rect 8562 4319 8878 4320
rect 5257 4314 5323 4317
rect 5901 4314 5967 4317
rect 18781 4314 18847 4317
rect 5257 4312 5967 4314
rect 5257 4256 5262 4312
rect 5318 4256 5906 4312
rect 5962 4256 5967 4312
rect 5257 4254 5967 4256
rect 5257 4251 5323 4254
rect 5901 4251 5967 4254
rect 9630 4312 18847 4314
rect 9630 4256 18786 4312
rect 18842 4256 18847 4312
rect 9630 4254 18847 4256
rect 2405 4178 2471 4181
rect 3969 4178 4035 4181
rect 9630 4178 9690 4254
rect 18781 4251 18847 4254
rect 2405 4176 2698 4178
rect 2405 4120 2410 4176
rect 2466 4120 2698 4176
rect 2405 4118 2698 4120
rect 2405 4115 2471 4118
rect 2638 4045 2698 4118
rect 3969 4176 9690 4178
rect 3969 4120 3974 4176
rect 4030 4120 9690 4176
rect 3969 4118 9690 4120
rect 13721 4178 13787 4181
rect 17309 4178 17375 4181
rect 13721 4176 17375 4178
rect 13721 4120 13726 4176
rect 13782 4120 17314 4176
rect 17370 4120 17375 4176
rect 13721 4118 17375 4120
rect 3969 4115 4035 4118
rect 13721 4115 13787 4118
rect 17309 4115 17375 4118
rect 2405 4042 2471 4045
rect 2405 4040 2514 4042
rect 2405 3984 2410 4040
rect 2466 3984 2514 4040
rect 2405 3979 2514 3984
rect 2638 4040 2747 4045
rect 2638 3984 2686 4040
rect 2742 3984 2747 4040
rect 2638 3982 2747 3984
rect 2681 3979 2747 3982
rect 4061 4042 4127 4045
rect 18965 4042 19031 4045
rect 4061 4040 19031 4042
rect 4061 3984 4066 4040
rect 4122 3984 18970 4040
rect 19026 3984 19031 4040
rect 4061 3982 19031 3984
rect 4061 3979 4127 3982
rect 18965 3979 19031 3982
rect 2454 3400 2514 3979
rect 2589 3906 2655 3909
rect 3141 3906 3207 3909
rect 2589 3904 3207 3906
rect 2589 3848 2594 3904
rect 2650 3848 3146 3904
rect 3202 3848 3207 3904
rect 2589 3846 3207 3848
rect 2589 3843 2655 3846
rect 3141 3843 3207 3846
rect 3325 3906 3391 3909
rect 4337 3906 4403 3909
rect 3325 3904 4403 3906
rect 3325 3848 3330 3904
rect 3386 3848 4342 3904
rect 4398 3848 4403 3904
rect 3325 3846 4403 3848
rect 3325 3843 3391 3846
rect 4337 3843 4403 3846
rect 9213 3906 9279 3909
rect 18045 3906 18111 3909
rect 9213 3904 18111 3906
rect 9213 3848 9218 3904
rect 9274 3848 18050 3904
rect 18106 3848 18111 3904
rect 9213 3846 18111 3848
rect 9213 3843 9279 3846
rect 18045 3843 18111 3846
rect 7562 3840 7878 3841
rect 7562 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7878 3840
rect 7562 3775 7878 3776
rect 2681 3770 2747 3773
rect 5441 3770 5507 3773
rect 2681 3768 5507 3770
rect 2681 3712 2686 3768
rect 2742 3712 5446 3768
rect 5502 3712 5507 3768
rect 2681 3710 5507 3712
rect 2681 3707 2747 3710
rect 5441 3707 5507 3710
rect 8201 3770 8267 3773
rect 12617 3770 12683 3773
rect 8201 3768 12683 3770
rect 8201 3712 8206 3768
rect 8262 3712 12622 3768
rect 12678 3712 12683 3768
rect 8201 3710 12683 3712
rect 8201 3707 8267 3710
rect 12617 3707 12683 3710
rect 13813 3770 13879 3773
rect 18321 3770 18387 3773
rect 13813 3768 18387 3770
rect 13813 3712 13818 3768
rect 13874 3712 18326 3768
rect 18382 3712 18387 3768
rect 13813 3710 18387 3712
rect 13813 3707 13879 3710
rect 18321 3707 18387 3710
rect 3141 3634 3207 3637
rect 6085 3634 6151 3637
rect 3141 3632 6151 3634
rect 3141 3576 3146 3632
rect 3202 3576 6090 3632
rect 6146 3576 6151 3632
rect 3141 3574 6151 3576
rect 3141 3571 3207 3574
rect 6085 3571 6151 3574
rect 7005 3634 7071 3637
rect 9765 3634 9831 3637
rect 7005 3632 9831 3634
rect 7005 3576 7010 3632
rect 7066 3576 9770 3632
rect 9826 3576 9831 3632
rect 7005 3574 9831 3576
rect 7005 3571 7071 3574
rect 9765 3571 9831 3574
rect 9949 3634 10015 3637
rect 12801 3634 12867 3637
rect 9949 3632 12867 3634
rect 9949 3576 9954 3632
rect 10010 3576 12806 3632
rect 12862 3576 12867 3632
rect 9949 3574 12867 3576
rect 9949 3571 10015 3574
rect 12801 3571 12867 3574
rect 7189 3498 7255 3501
rect 9213 3498 9279 3501
rect 11513 3498 11579 3501
rect 7189 3496 9138 3498
rect 7189 3440 7194 3496
rect 7250 3440 9138 3496
rect 7189 3438 9138 3440
rect 7189 3435 7255 3438
rect 5533 3362 5599 3365
rect 7925 3362 7991 3365
rect 5533 3360 7991 3362
rect 5533 3304 5538 3360
rect 5594 3304 7930 3360
rect 7986 3304 7991 3360
rect 5533 3302 7991 3304
rect 9078 3362 9138 3438
rect 9213 3496 11579 3498
rect 9213 3440 9218 3496
rect 9274 3440 11518 3496
rect 11574 3440 11579 3496
rect 9213 3438 11579 3440
rect 9213 3435 9279 3438
rect 11513 3435 11579 3438
rect 11053 3362 11119 3365
rect 9078 3360 11119 3362
rect 9078 3304 11058 3360
rect 11114 3304 11119 3360
rect 9078 3302 11119 3304
rect 5533 3299 5599 3302
rect 7925 3299 7991 3302
rect 11053 3299 11119 3302
rect 11697 3362 11763 3365
rect 12985 3362 13051 3365
rect 11697 3360 13051 3362
rect 11697 3304 11702 3360
rect 11758 3304 12990 3360
rect 13046 3304 13051 3360
rect 11697 3302 13051 3304
rect 11697 3299 11763 3302
rect 12985 3299 13051 3302
rect 3562 3296 3878 3297
rect 3562 3232 3568 3296
rect 3632 3232 3648 3296
rect 3712 3232 3728 3296
rect 3792 3232 3808 3296
rect 3872 3232 3878 3296
rect 3562 3231 3878 3232
rect 8562 3296 8878 3297
rect 8562 3232 8568 3296
rect 8632 3232 8648 3296
rect 8712 3232 8728 3296
rect 8792 3232 8808 3296
rect 8872 3232 8878 3296
rect 8562 3231 8878 3232
rect 6085 3226 6151 3229
rect 8293 3226 8359 3229
rect 6085 3224 8359 3226
rect 6085 3168 6090 3224
rect 6146 3168 8298 3224
rect 8354 3168 8359 3224
rect 6085 3166 8359 3168
rect 6085 3163 6151 3166
rect 8293 3163 8359 3166
rect 9121 3226 9187 3229
rect 12249 3226 12315 3229
rect 9121 3224 12315 3226
rect 9121 3168 9126 3224
rect 9182 3168 12254 3224
rect 12310 3168 12315 3224
rect 9121 3166 12315 3168
rect 9121 3163 9187 3166
rect 12249 3163 12315 3166
rect 5349 3090 5415 3093
rect 19057 3090 19123 3093
rect 5349 3088 19123 3090
rect 5349 3032 5354 3088
rect 5410 3032 19062 3088
rect 19118 3032 19123 3088
rect 5349 3030 19123 3032
rect 5349 3027 5415 3030
rect 19057 3027 19123 3030
rect 6545 2954 6611 2957
rect 9029 2954 9095 2957
rect 6545 2952 9095 2954
rect 6545 2896 6550 2952
rect 6606 2896 9034 2952
rect 9090 2896 9095 2952
rect 6545 2894 9095 2896
rect 6545 2891 6611 2894
rect 9029 2891 9095 2894
rect 9213 2954 9279 2957
rect 10869 2954 10935 2957
rect 9213 2952 10935 2954
rect 9213 2896 9218 2952
rect 9274 2896 10874 2952
rect 10930 2896 10935 2952
rect 9213 2894 10935 2896
rect 9213 2891 9279 2894
rect 10869 2891 10935 2894
rect 8753 2818 8819 2821
rect 12341 2818 12407 2821
rect 8753 2816 12407 2818
rect 8753 2760 8758 2816
rect 8814 2760 12346 2816
rect 12402 2760 12407 2816
rect 8753 2758 12407 2760
rect 8753 2755 8819 2758
rect 12341 2755 12407 2758
rect 7562 2752 7878 2753
rect 7562 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7878 2752
rect 7562 2687 7878 2688
rect 2497 2682 2563 2685
rect 5901 2682 5967 2685
rect 2497 2680 5967 2682
rect 2497 2624 2502 2680
rect 2558 2624 5906 2680
rect 5962 2624 5967 2680
rect 2497 2622 5967 2624
rect 2497 2619 2563 2622
rect 5901 2619 5967 2622
rect 8334 2620 8340 2684
rect 8404 2682 8410 2684
rect 9213 2682 9279 2685
rect 8404 2680 9279 2682
rect 8404 2624 9218 2680
rect 9274 2624 9279 2680
rect 8404 2622 9279 2624
rect 8404 2620 8410 2622
rect 9213 2619 9279 2622
rect 2681 2546 2747 2549
rect 5625 2546 5691 2549
rect 2681 2544 5691 2546
rect 2681 2488 2686 2544
rect 2742 2488 5630 2544
rect 5686 2488 5691 2544
rect 2681 2486 5691 2488
rect 2681 2483 2747 2486
rect 5625 2483 5691 2486
rect 6637 2546 6703 2549
rect 18045 2546 18111 2549
rect 6637 2544 18111 2546
rect 6637 2488 6642 2544
rect 6698 2488 18050 2544
rect 18106 2488 18111 2544
rect 6637 2486 18111 2488
rect 6637 2483 6703 2486
rect 18045 2483 18111 2486
rect 5441 2410 5507 2413
rect 8753 2410 8819 2413
rect 5441 2408 8819 2410
rect 5441 2352 5446 2408
rect 5502 2352 8758 2408
rect 8814 2352 8819 2408
rect 5441 2350 8819 2352
rect 5441 2347 5507 2350
rect 8753 2347 8819 2350
rect 8937 2410 9003 2413
rect 16849 2410 16915 2413
rect 8937 2408 16915 2410
rect 8937 2352 8942 2408
rect 8998 2352 16854 2408
rect 16910 2352 16915 2408
rect 8937 2350 16915 2352
rect 8937 2347 9003 2350
rect 16849 2347 16915 2350
rect 4705 2274 4771 2277
rect 8385 2274 8451 2277
rect 4705 2272 8451 2274
rect 4705 2216 4710 2272
rect 4766 2216 8390 2272
rect 8446 2216 8451 2272
rect 4705 2214 8451 2216
rect 4705 2211 4771 2214
rect 8385 2211 8451 2214
rect 9029 2274 9095 2277
rect 12065 2274 12131 2277
rect 9029 2272 12131 2274
rect 9029 2216 9034 2272
rect 9090 2216 12070 2272
rect 12126 2216 12131 2272
rect 9029 2214 12131 2216
rect 9029 2211 9095 2214
rect 12065 2211 12131 2214
rect 3562 2208 3878 2209
rect 3562 2144 3568 2208
rect 3632 2144 3648 2208
rect 3712 2144 3728 2208
rect 3792 2144 3808 2208
rect 3872 2144 3878 2208
rect 3562 2143 3878 2144
rect 8562 2208 8878 2209
rect 8562 2144 8568 2208
rect 8632 2144 8648 2208
rect 8712 2144 8728 2208
rect 8792 2144 8808 2208
rect 8872 2144 8878 2208
rect 8562 2143 8878 2144
rect 6729 2138 6795 2141
rect 8150 2138 8156 2140
rect 6729 2136 8156 2138
rect 6729 2080 6734 2136
rect 6790 2080 8156 2136
rect 6729 2078 8156 2080
rect 6729 2075 6795 2078
rect 8150 2076 8156 2078
rect 8220 2076 8226 2140
rect 9305 2138 9371 2141
rect 9581 2138 9647 2141
rect 18413 2138 18479 2141
rect 9305 2136 18479 2138
rect 9305 2080 9310 2136
rect 9366 2080 9586 2136
rect 9642 2080 18418 2136
rect 18474 2080 18479 2136
rect 9305 2078 18479 2080
rect 9305 2075 9371 2078
rect 9581 2075 9647 2078
rect 18413 2075 18479 2078
rect 5625 2002 5691 2005
rect 13813 2002 13879 2005
rect 5625 2000 13879 2002
rect 5625 1944 5630 2000
rect 5686 1944 13818 2000
rect 13874 1944 13879 2000
rect 5625 1942 13879 1944
rect 5625 1939 5691 1942
rect 13813 1939 13879 1942
rect 7465 1866 7531 1869
rect 11237 1866 11303 1869
rect 7465 1864 11303 1866
rect 7465 1808 7470 1864
rect 7526 1808 11242 1864
rect 11298 1808 11303 1864
rect 7465 1806 11303 1808
rect 7465 1803 7531 1806
rect 11237 1803 11303 1806
rect 2865 1730 2931 1733
rect 5993 1730 6059 1733
rect 2865 1728 6059 1730
rect 2865 1672 2870 1728
rect 2926 1672 5998 1728
rect 6054 1672 6059 1728
rect 2865 1670 6059 1672
rect 2865 1667 2931 1670
rect 5993 1667 6059 1670
rect 8385 1730 8451 1733
rect 11697 1730 11763 1733
rect 8385 1728 11763 1730
rect 8385 1672 8390 1728
rect 8446 1672 11702 1728
rect 11758 1672 11763 1728
rect 8385 1670 11763 1672
rect 8385 1667 8451 1670
rect 11697 1667 11763 1670
rect 7562 1664 7878 1665
rect 7562 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7878 1664
rect 7562 1599 7878 1600
rect 289 1594 355 1597
rect 1853 1594 1919 1597
rect 289 1592 1919 1594
rect 289 1536 294 1592
rect 350 1536 1858 1592
rect 1914 1536 1919 1592
rect 289 1534 1919 1536
rect 289 1531 355 1534
rect 1853 1531 1919 1534
rect 2313 1594 2379 1597
rect 4153 1594 4219 1597
rect 2313 1592 4219 1594
rect 2313 1536 2318 1592
rect 2374 1536 4158 1592
rect 4214 1536 4219 1592
rect 2313 1534 4219 1536
rect 2313 1531 2379 1534
rect 4153 1531 4219 1534
rect 8150 1532 8156 1596
rect 8220 1594 8226 1596
rect 16941 1594 17007 1597
rect 8220 1592 17007 1594
rect 8220 1536 16946 1592
rect 17002 1536 17007 1592
rect 8220 1534 17007 1536
rect 8220 1532 8226 1534
rect 16941 1531 17007 1534
rect 933 1458 999 1461
rect 2773 1458 2839 1461
rect 933 1456 2839 1458
rect 933 1400 938 1456
rect 994 1400 2778 1456
rect 2834 1400 2839 1456
rect 933 1398 2839 1400
rect 933 1395 999 1398
rect 2773 1395 2839 1398
rect 6177 1458 6243 1461
rect 15101 1458 15167 1461
rect 6177 1456 15167 1458
rect 6177 1400 6182 1456
rect 6238 1400 15106 1456
rect 15162 1400 15167 1456
rect 6177 1398 15167 1400
rect 6177 1395 6243 1398
rect 15101 1395 15167 1398
rect 1117 1322 1183 1325
rect 3601 1322 3667 1325
rect 1117 1320 3667 1322
rect 1117 1264 1122 1320
rect 1178 1264 3606 1320
rect 3662 1264 3667 1320
rect 1117 1262 3667 1264
rect 1117 1259 1183 1262
rect 3601 1259 3667 1262
rect 4061 1322 4127 1325
rect 7373 1322 7439 1325
rect 4061 1320 7439 1322
rect 4061 1264 4066 1320
rect 4122 1264 7378 1320
rect 7434 1264 7439 1320
rect 4061 1262 7439 1264
rect 4061 1259 4127 1262
rect 7373 1259 7439 1262
rect 8201 1322 8267 1325
rect 18505 1322 18571 1325
rect 8201 1320 18571 1322
rect 8201 1264 8206 1320
rect 8262 1264 18510 1320
rect 18566 1264 18571 1320
rect 8201 1262 18571 1264
rect 8201 1259 8267 1262
rect 18505 1259 18571 1262
rect 565 1186 631 1189
rect 2865 1186 2931 1189
rect 565 1184 2931 1186
rect 565 1128 570 1184
rect 626 1128 2870 1184
rect 2926 1128 2931 1184
rect 565 1126 2931 1128
rect 565 1123 631 1126
rect 2865 1123 2931 1126
rect 3562 1120 3878 1121
rect 3562 1056 3568 1120
rect 3632 1056 3648 1120
rect 3712 1056 3728 1120
rect 3792 1056 3808 1120
rect 3872 1056 3878 1120
rect 3562 1055 3878 1056
rect 8562 1120 8878 1121
rect 8562 1056 8568 1120
rect 8632 1056 8648 1120
rect 8712 1056 8728 1120
rect 8792 1056 8808 1120
rect 8872 1056 8878 1120
rect 8562 1055 8878 1056
rect 5993 1050 6059 1053
rect 3972 1048 6059 1050
rect 3972 992 5998 1048
rect 6054 992 6059 1048
rect 3972 990 6059 992
rect 1025 914 1091 917
rect 3972 914 4032 990
rect 5993 987 6059 990
rect 1025 912 4032 914
rect 1025 856 1030 912
rect 1086 856 4032 912
rect 1025 854 4032 856
rect 4889 914 4955 917
rect 14273 914 14339 917
rect 4889 912 14339 914
rect 4889 856 4894 912
rect 4950 856 14278 912
rect 14334 856 14339 912
rect 4889 854 14339 856
rect 1025 851 1091 854
rect 4889 851 4955 854
rect 14273 851 14339 854
rect 4337 778 4403 781
rect 17769 778 17835 781
rect 4337 776 17835 778
rect 4337 720 4342 776
rect 4398 720 17774 776
rect 17830 720 17835 776
rect 4337 718 17835 720
rect 4337 715 4403 718
rect 17769 715 17835 718
rect 4153 642 4219 645
rect 8109 642 8175 645
rect 4153 640 8175 642
rect 4153 584 4158 640
rect 4214 584 8114 640
rect 8170 584 8175 640
rect 4153 582 8175 584
rect 4153 579 4219 582
rect 8109 579 8175 582
rect 8293 642 8359 645
rect 17861 642 17927 645
rect 8293 640 17927 642
rect 8293 584 8298 640
rect 8354 584 17866 640
rect 17922 584 17927 640
rect 8293 582 17927 584
rect 8293 579 8359 582
rect 17861 579 17927 582
rect 9121 506 9187 509
rect 18597 506 18663 509
rect 9121 504 18663 506
rect 9121 448 9126 504
rect 9182 448 18602 504
rect 18658 448 18663 504
rect 9121 446 18663 448
rect 9121 443 9187 446
rect 18597 443 18663 446
rect 6729 370 6795 373
rect 13905 370 13971 373
rect 6729 368 13971 370
rect 6729 312 6734 368
rect 6790 312 13910 368
rect 13966 312 13971 368
rect 6729 310 13971 312
rect 6729 307 6795 310
rect 13905 307 13971 310
rect 8109 234 8175 237
rect 14089 234 14155 237
rect 8109 232 14155 234
rect 8109 176 8114 232
rect 8170 176 14094 232
rect 14150 176 14155 232
rect 8109 174 14155 176
rect 8109 171 8175 174
rect 14089 171 14155 174
<< via3 >>
rect 2568 15804 2632 15808
rect 2568 15748 2572 15804
rect 2572 15748 2628 15804
rect 2628 15748 2632 15804
rect 2568 15744 2632 15748
rect 2648 15804 2712 15808
rect 2648 15748 2652 15804
rect 2652 15748 2708 15804
rect 2708 15748 2712 15804
rect 2648 15744 2712 15748
rect 2728 15804 2792 15808
rect 2728 15748 2732 15804
rect 2732 15748 2788 15804
rect 2788 15748 2792 15804
rect 2728 15744 2792 15748
rect 2808 15804 2872 15808
rect 2808 15748 2812 15804
rect 2812 15748 2868 15804
rect 2868 15748 2872 15804
rect 2808 15744 2872 15748
rect 7568 15804 7632 15808
rect 7568 15748 7572 15804
rect 7572 15748 7628 15804
rect 7628 15748 7632 15804
rect 7568 15744 7632 15748
rect 7648 15804 7712 15808
rect 7648 15748 7652 15804
rect 7652 15748 7708 15804
rect 7708 15748 7712 15804
rect 7648 15744 7712 15748
rect 7728 15804 7792 15808
rect 7728 15748 7732 15804
rect 7732 15748 7788 15804
rect 7788 15748 7792 15804
rect 7728 15744 7792 15748
rect 7808 15804 7872 15808
rect 7808 15748 7812 15804
rect 7812 15748 7868 15804
rect 7868 15748 7872 15804
rect 7808 15744 7872 15748
rect 3568 15260 3632 15264
rect 3568 15204 3572 15260
rect 3572 15204 3628 15260
rect 3628 15204 3632 15260
rect 3568 15200 3632 15204
rect 3648 15260 3712 15264
rect 3648 15204 3652 15260
rect 3652 15204 3708 15260
rect 3708 15204 3712 15260
rect 3648 15200 3712 15204
rect 3728 15260 3792 15264
rect 3728 15204 3732 15260
rect 3732 15204 3788 15260
rect 3788 15204 3792 15260
rect 3728 15200 3792 15204
rect 3808 15260 3872 15264
rect 3808 15204 3812 15260
rect 3812 15204 3868 15260
rect 3868 15204 3872 15260
rect 3808 15200 3872 15204
rect 8568 15260 8632 15264
rect 8568 15204 8572 15260
rect 8572 15204 8628 15260
rect 8628 15204 8632 15260
rect 8568 15200 8632 15204
rect 8648 15260 8712 15264
rect 8648 15204 8652 15260
rect 8652 15204 8708 15260
rect 8708 15204 8712 15260
rect 8648 15200 8712 15204
rect 8728 15260 8792 15264
rect 8728 15204 8732 15260
rect 8732 15204 8788 15260
rect 8788 15204 8792 15260
rect 8728 15200 8792 15204
rect 8808 15260 8872 15264
rect 8808 15204 8812 15260
rect 8812 15204 8868 15260
rect 8868 15204 8872 15260
rect 8808 15200 8872 15204
rect 2568 14716 2632 14720
rect 2568 14660 2572 14716
rect 2572 14660 2628 14716
rect 2628 14660 2632 14716
rect 2568 14656 2632 14660
rect 2648 14716 2712 14720
rect 2648 14660 2652 14716
rect 2652 14660 2708 14716
rect 2708 14660 2712 14716
rect 2648 14656 2712 14660
rect 2728 14716 2792 14720
rect 2728 14660 2732 14716
rect 2732 14660 2788 14716
rect 2788 14660 2792 14716
rect 2728 14656 2792 14660
rect 2808 14716 2872 14720
rect 2808 14660 2812 14716
rect 2812 14660 2868 14716
rect 2868 14660 2872 14716
rect 2808 14656 2872 14660
rect 7568 14716 7632 14720
rect 7568 14660 7572 14716
rect 7572 14660 7628 14716
rect 7628 14660 7632 14716
rect 7568 14656 7632 14660
rect 7648 14716 7712 14720
rect 7648 14660 7652 14716
rect 7652 14660 7708 14716
rect 7708 14660 7712 14716
rect 7648 14656 7712 14660
rect 7728 14716 7792 14720
rect 7728 14660 7732 14716
rect 7732 14660 7788 14716
rect 7788 14660 7792 14716
rect 7728 14656 7792 14660
rect 7808 14716 7872 14720
rect 7808 14660 7812 14716
rect 7812 14660 7868 14716
rect 7868 14660 7872 14716
rect 7808 14656 7872 14660
rect 3568 14172 3632 14176
rect 3568 14116 3572 14172
rect 3572 14116 3628 14172
rect 3628 14116 3632 14172
rect 3568 14112 3632 14116
rect 3648 14172 3712 14176
rect 3648 14116 3652 14172
rect 3652 14116 3708 14172
rect 3708 14116 3712 14172
rect 3648 14112 3712 14116
rect 3728 14172 3792 14176
rect 3728 14116 3732 14172
rect 3732 14116 3788 14172
rect 3788 14116 3792 14172
rect 3728 14112 3792 14116
rect 3808 14172 3872 14176
rect 3808 14116 3812 14172
rect 3812 14116 3868 14172
rect 3868 14116 3872 14172
rect 3808 14112 3872 14116
rect 8568 14172 8632 14176
rect 8568 14116 8572 14172
rect 8572 14116 8628 14172
rect 8628 14116 8632 14172
rect 8568 14112 8632 14116
rect 8648 14172 8712 14176
rect 8648 14116 8652 14172
rect 8652 14116 8708 14172
rect 8708 14116 8712 14172
rect 8648 14112 8712 14116
rect 8728 14172 8792 14176
rect 8728 14116 8732 14172
rect 8732 14116 8788 14172
rect 8788 14116 8792 14172
rect 8728 14112 8792 14116
rect 8808 14172 8872 14176
rect 8808 14116 8812 14172
rect 8812 14116 8868 14172
rect 8868 14116 8872 14172
rect 8808 14112 8872 14116
rect 7236 13772 7300 13836
rect 2568 13628 2632 13632
rect 2568 13572 2572 13628
rect 2572 13572 2628 13628
rect 2628 13572 2632 13628
rect 2568 13568 2632 13572
rect 2648 13628 2712 13632
rect 2648 13572 2652 13628
rect 2652 13572 2708 13628
rect 2708 13572 2712 13628
rect 2648 13568 2712 13572
rect 2728 13628 2792 13632
rect 2728 13572 2732 13628
rect 2732 13572 2788 13628
rect 2788 13572 2792 13628
rect 2728 13568 2792 13572
rect 2808 13628 2872 13632
rect 2808 13572 2812 13628
rect 2812 13572 2868 13628
rect 2868 13572 2872 13628
rect 2808 13568 2872 13572
rect 7568 13628 7632 13632
rect 7568 13572 7572 13628
rect 7572 13572 7628 13628
rect 7628 13572 7632 13628
rect 7568 13568 7632 13572
rect 7648 13628 7712 13632
rect 7648 13572 7652 13628
rect 7652 13572 7708 13628
rect 7708 13572 7712 13628
rect 7648 13568 7712 13572
rect 7728 13628 7792 13632
rect 7728 13572 7732 13628
rect 7732 13572 7788 13628
rect 7788 13572 7792 13628
rect 7728 13568 7792 13572
rect 7808 13628 7872 13632
rect 7808 13572 7812 13628
rect 7812 13572 7868 13628
rect 7868 13572 7872 13628
rect 7808 13568 7872 13572
rect 3568 13084 3632 13088
rect 3568 13028 3572 13084
rect 3572 13028 3628 13084
rect 3628 13028 3632 13084
rect 3568 13024 3632 13028
rect 3648 13084 3712 13088
rect 3648 13028 3652 13084
rect 3652 13028 3708 13084
rect 3708 13028 3712 13084
rect 3648 13024 3712 13028
rect 3728 13084 3792 13088
rect 3728 13028 3732 13084
rect 3732 13028 3788 13084
rect 3788 13028 3792 13084
rect 3728 13024 3792 13028
rect 3808 13084 3872 13088
rect 3808 13028 3812 13084
rect 3812 13028 3868 13084
rect 3868 13028 3872 13084
rect 3808 13024 3872 13028
rect 8568 13084 8632 13088
rect 8568 13028 8572 13084
rect 8572 13028 8628 13084
rect 8628 13028 8632 13084
rect 8568 13024 8632 13028
rect 8648 13084 8712 13088
rect 8648 13028 8652 13084
rect 8652 13028 8708 13084
rect 8708 13028 8712 13084
rect 8648 13024 8712 13028
rect 8728 13084 8792 13088
rect 8728 13028 8732 13084
rect 8732 13028 8788 13084
rect 8788 13028 8792 13084
rect 8728 13024 8792 13028
rect 8808 13084 8872 13088
rect 8808 13028 8812 13084
rect 8812 13028 8868 13084
rect 8868 13028 8872 13084
rect 8808 13024 8872 13028
rect 2568 12540 2632 12544
rect 2568 12484 2572 12540
rect 2572 12484 2628 12540
rect 2628 12484 2632 12540
rect 2568 12480 2632 12484
rect 2648 12540 2712 12544
rect 2648 12484 2652 12540
rect 2652 12484 2708 12540
rect 2708 12484 2712 12540
rect 2648 12480 2712 12484
rect 2728 12540 2792 12544
rect 2728 12484 2732 12540
rect 2732 12484 2788 12540
rect 2788 12484 2792 12540
rect 2728 12480 2792 12484
rect 2808 12540 2872 12544
rect 2808 12484 2812 12540
rect 2812 12484 2868 12540
rect 2868 12484 2872 12540
rect 2808 12480 2872 12484
rect 7568 12540 7632 12544
rect 7568 12484 7572 12540
rect 7572 12484 7628 12540
rect 7628 12484 7632 12540
rect 7568 12480 7632 12484
rect 7648 12540 7712 12544
rect 7648 12484 7652 12540
rect 7652 12484 7708 12540
rect 7708 12484 7712 12540
rect 7648 12480 7712 12484
rect 7728 12540 7792 12544
rect 7728 12484 7732 12540
rect 7732 12484 7788 12540
rect 7788 12484 7792 12540
rect 7728 12480 7792 12484
rect 7808 12540 7872 12544
rect 7808 12484 7812 12540
rect 7812 12484 7868 12540
rect 7868 12484 7872 12540
rect 7808 12480 7872 12484
rect 1348 12276 1412 12340
rect 1348 12064 1412 12068
rect 1348 12008 1362 12064
rect 1362 12008 1412 12064
rect 1348 12004 1412 12008
rect 3568 11996 3632 12000
rect 3568 11940 3572 11996
rect 3572 11940 3628 11996
rect 3628 11940 3632 11996
rect 3568 11936 3632 11940
rect 3648 11996 3712 12000
rect 3648 11940 3652 11996
rect 3652 11940 3708 11996
rect 3708 11940 3712 11996
rect 3648 11936 3712 11940
rect 3728 11996 3792 12000
rect 3728 11940 3732 11996
rect 3732 11940 3788 11996
rect 3788 11940 3792 11996
rect 3728 11936 3792 11940
rect 3808 11996 3872 12000
rect 3808 11940 3812 11996
rect 3812 11940 3868 11996
rect 3868 11940 3872 11996
rect 3808 11936 3872 11940
rect 8568 11996 8632 12000
rect 8568 11940 8572 11996
rect 8572 11940 8628 11996
rect 8628 11940 8632 11996
rect 8568 11936 8632 11940
rect 8648 11996 8712 12000
rect 8648 11940 8652 11996
rect 8652 11940 8708 11996
rect 8708 11940 8712 11996
rect 8648 11936 8712 11940
rect 8728 11996 8792 12000
rect 8728 11940 8732 11996
rect 8732 11940 8788 11996
rect 8788 11940 8792 11996
rect 8728 11936 8792 11940
rect 8808 11996 8872 12000
rect 8808 11940 8812 11996
rect 8812 11940 8868 11996
rect 8868 11940 8872 11996
rect 8808 11936 8872 11940
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 7568 11452 7632 11456
rect 7568 11396 7572 11452
rect 7572 11396 7628 11452
rect 7628 11396 7632 11452
rect 7568 11392 7632 11396
rect 7648 11452 7712 11456
rect 7648 11396 7652 11452
rect 7652 11396 7708 11452
rect 7708 11396 7712 11452
rect 7648 11392 7712 11396
rect 7728 11452 7792 11456
rect 7728 11396 7732 11452
rect 7732 11396 7788 11452
rect 7788 11396 7792 11452
rect 7728 11392 7792 11396
rect 7808 11452 7872 11456
rect 7808 11396 7812 11452
rect 7812 11396 7868 11452
rect 7868 11396 7872 11452
rect 7808 11392 7872 11396
rect 3568 10908 3632 10912
rect 3568 10852 3572 10908
rect 3572 10852 3628 10908
rect 3628 10852 3632 10908
rect 3568 10848 3632 10852
rect 3648 10908 3712 10912
rect 3648 10852 3652 10908
rect 3652 10852 3708 10908
rect 3708 10852 3712 10908
rect 3648 10848 3712 10852
rect 3728 10908 3792 10912
rect 3728 10852 3732 10908
rect 3732 10852 3788 10908
rect 3788 10852 3792 10908
rect 3728 10848 3792 10852
rect 3808 10908 3872 10912
rect 3808 10852 3812 10908
rect 3812 10852 3868 10908
rect 3868 10852 3872 10908
rect 3808 10848 3872 10852
rect 8568 10908 8632 10912
rect 8568 10852 8572 10908
rect 8572 10852 8628 10908
rect 8628 10852 8632 10908
rect 8568 10848 8632 10852
rect 8648 10908 8712 10912
rect 8648 10852 8652 10908
rect 8652 10852 8708 10908
rect 8708 10852 8712 10908
rect 8648 10848 8712 10852
rect 8728 10908 8792 10912
rect 8728 10852 8732 10908
rect 8732 10852 8788 10908
rect 8788 10852 8792 10908
rect 8728 10848 8792 10852
rect 8808 10908 8872 10912
rect 8808 10852 8812 10908
rect 8812 10852 8868 10908
rect 8868 10852 8872 10908
rect 8808 10848 8872 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 7568 10364 7632 10368
rect 7568 10308 7572 10364
rect 7572 10308 7628 10364
rect 7628 10308 7632 10364
rect 7568 10304 7632 10308
rect 7648 10364 7712 10368
rect 7648 10308 7652 10364
rect 7652 10308 7708 10364
rect 7708 10308 7712 10364
rect 7648 10304 7712 10308
rect 7728 10364 7792 10368
rect 7728 10308 7732 10364
rect 7732 10308 7788 10364
rect 7788 10308 7792 10364
rect 7728 10304 7792 10308
rect 7808 10364 7872 10368
rect 7808 10308 7812 10364
rect 7812 10308 7868 10364
rect 7868 10308 7872 10364
rect 7808 10304 7872 10308
rect 3568 9820 3632 9824
rect 3568 9764 3572 9820
rect 3572 9764 3628 9820
rect 3628 9764 3632 9820
rect 3568 9760 3632 9764
rect 3648 9820 3712 9824
rect 3648 9764 3652 9820
rect 3652 9764 3708 9820
rect 3708 9764 3712 9820
rect 3648 9760 3712 9764
rect 3728 9820 3792 9824
rect 3728 9764 3732 9820
rect 3732 9764 3788 9820
rect 3788 9764 3792 9820
rect 3728 9760 3792 9764
rect 3808 9820 3872 9824
rect 3808 9764 3812 9820
rect 3812 9764 3868 9820
rect 3868 9764 3872 9820
rect 3808 9760 3872 9764
rect 8568 9820 8632 9824
rect 8568 9764 8572 9820
rect 8572 9764 8628 9820
rect 8628 9764 8632 9820
rect 8568 9760 8632 9764
rect 8648 9820 8712 9824
rect 8648 9764 8652 9820
rect 8652 9764 8708 9820
rect 8708 9764 8712 9820
rect 8648 9760 8712 9764
rect 8728 9820 8792 9824
rect 8728 9764 8732 9820
rect 8732 9764 8788 9820
rect 8788 9764 8792 9820
rect 8728 9760 8792 9764
rect 8808 9820 8872 9824
rect 8808 9764 8812 9820
rect 8812 9764 8868 9820
rect 8868 9764 8872 9820
rect 8808 9760 8872 9764
rect 7236 9284 7300 9348
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 7568 9276 7632 9280
rect 7568 9220 7572 9276
rect 7572 9220 7628 9276
rect 7628 9220 7632 9276
rect 7568 9216 7632 9220
rect 7648 9276 7712 9280
rect 7648 9220 7652 9276
rect 7652 9220 7708 9276
rect 7708 9220 7712 9276
rect 7648 9216 7712 9220
rect 7728 9276 7792 9280
rect 7728 9220 7732 9276
rect 7732 9220 7788 9276
rect 7788 9220 7792 9276
rect 7728 9216 7792 9220
rect 7808 9276 7872 9280
rect 7808 9220 7812 9276
rect 7812 9220 7868 9276
rect 7868 9220 7872 9276
rect 7808 9216 7872 9220
rect 8340 8876 8404 8940
rect 3568 8732 3632 8736
rect 3568 8676 3572 8732
rect 3572 8676 3628 8732
rect 3628 8676 3632 8732
rect 3568 8672 3632 8676
rect 3648 8732 3712 8736
rect 3648 8676 3652 8732
rect 3652 8676 3708 8732
rect 3708 8676 3712 8732
rect 3648 8672 3712 8676
rect 3728 8732 3792 8736
rect 3728 8676 3732 8732
rect 3732 8676 3788 8732
rect 3788 8676 3792 8732
rect 3728 8672 3792 8676
rect 3808 8732 3872 8736
rect 3808 8676 3812 8732
rect 3812 8676 3868 8732
rect 3868 8676 3872 8732
rect 3808 8672 3872 8676
rect 8568 8732 8632 8736
rect 8568 8676 8572 8732
rect 8572 8676 8628 8732
rect 8628 8676 8632 8732
rect 8568 8672 8632 8676
rect 8648 8732 8712 8736
rect 8648 8676 8652 8732
rect 8652 8676 8708 8732
rect 8708 8676 8712 8732
rect 8648 8672 8712 8676
rect 8728 8732 8792 8736
rect 8728 8676 8732 8732
rect 8732 8676 8788 8732
rect 8788 8676 8792 8732
rect 8728 8672 8792 8676
rect 8808 8732 8872 8736
rect 8808 8676 8812 8732
rect 8812 8676 8868 8732
rect 8868 8676 8872 8732
rect 8808 8672 8872 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 7568 8188 7632 8192
rect 7568 8132 7572 8188
rect 7572 8132 7628 8188
rect 7628 8132 7632 8188
rect 7568 8128 7632 8132
rect 7648 8188 7712 8192
rect 7648 8132 7652 8188
rect 7652 8132 7708 8188
rect 7708 8132 7712 8188
rect 7648 8128 7712 8132
rect 7728 8188 7792 8192
rect 7728 8132 7732 8188
rect 7732 8132 7788 8188
rect 7788 8132 7792 8188
rect 7728 8128 7792 8132
rect 7808 8188 7872 8192
rect 7808 8132 7812 8188
rect 7812 8132 7868 8188
rect 7868 8132 7872 8188
rect 7808 8128 7872 8132
rect 3568 7644 3632 7648
rect 3568 7588 3572 7644
rect 3572 7588 3628 7644
rect 3628 7588 3632 7644
rect 3568 7584 3632 7588
rect 3648 7644 3712 7648
rect 3648 7588 3652 7644
rect 3652 7588 3708 7644
rect 3708 7588 3712 7644
rect 3648 7584 3712 7588
rect 3728 7644 3792 7648
rect 3728 7588 3732 7644
rect 3732 7588 3788 7644
rect 3788 7588 3792 7644
rect 3728 7584 3792 7588
rect 3808 7644 3872 7648
rect 3808 7588 3812 7644
rect 3812 7588 3868 7644
rect 3868 7588 3872 7644
rect 3808 7584 3872 7588
rect 8568 7644 8632 7648
rect 8568 7588 8572 7644
rect 8572 7588 8628 7644
rect 8628 7588 8632 7644
rect 8568 7584 8632 7588
rect 8648 7644 8712 7648
rect 8648 7588 8652 7644
rect 8652 7588 8708 7644
rect 8708 7588 8712 7644
rect 8648 7584 8712 7588
rect 8728 7644 8792 7648
rect 8728 7588 8732 7644
rect 8732 7588 8788 7644
rect 8788 7588 8792 7644
rect 8728 7584 8792 7588
rect 8808 7644 8872 7648
rect 8808 7588 8812 7644
rect 8812 7588 8868 7644
rect 8868 7588 8872 7644
rect 8808 7584 8872 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 7568 7100 7632 7104
rect 7568 7044 7572 7100
rect 7572 7044 7628 7100
rect 7628 7044 7632 7100
rect 7568 7040 7632 7044
rect 7648 7100 7712 7104
rect 7648 7044 7652 7100
rect 7652 7044 7708 7100
rect 7708 7044 7712 7100
rect 7648 7040 7712 7044
rect 7728 7100 7792 7104
rect 7728 7044 7732 7100
rect 7732 7044 7788 7100
rect 7788 7044 7792 7100
rect 7728 7040 7792 7044
rect 7808 7100 7872 7104
rect 7808 7044 7812 7100
rect 7812 7044 7868 7100
rect 7868 7044 7872 7100
rect 7808 7040 7872 7044
rect 3568 6556 3632 6560
rect 3568 6500 3572 6556
rect 3572 6500 3628 6556
rect 3628 6500 3632 6556
rect 3568 6496 3632 6500
rect 3648 6556 3712 6560
rect 3648 6500 3652 6556
rect 3652 6500 3708 6556
rect 3708 6500 3712 6556
rect 3648 6496 3712 6500
rect 3728 6556 3792 6560
rect 3728 6500 3732 6556
rect 3732 6500 3788 6556
rect 3788 6500 3792 6556
rect 3728 6496 3792 6500
rect 3808 6556 3872 6560
rect 3808 6500 3812 6556
rect 3812 6500 3868 6556
rect 3868 6500 3872 6556
rect 3808 6496 3872 6500
rect 8568 6556 8632 6560
rect 8568 6500 8572 6556
rect 8572 6500 8628 6556
rect 8628 6500 8632 6556
rect 8568 6496 8632 6500
rect 8648 6556 8712 6560
rect 8648 6500 8652 6556
rect 8652 6500 8708 6556
rect 8708 6500 8712 6556
rect 8648 6496 8712 6500
rect 8728 6556 8792 6560
rect 8728 6500 8732 6556
rect 8732 6500 8788 6556
rect 8788 6500 8792 6556
rect 8728 6496 8792 6500
rect 8808 6556 8872 6560
rect 8808 6500 8812 6556
rect 8812 6500 8868 6556
rect 8868 6500 8872 6556
rect 8808 6496 8872 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 7568 6012 7632 6016
rect 7568 5956 7572 6012
rect 7572 5956 7628 6012
rect 7628 5956 7632 6012
rect 7568 5952 7632 5956
rect 7648 6012 7712 6016
rect 7648 5956 7652 6012
rect 7652 5956 7708 6012
rect 7708 5956 7712 6012
rect 7648 5952 7712 5956
rect 7728 6012 7792 6016
rect 7728 5956 7732 6012
rect 7732 5956 7788 6012
rect 7788 5956 7792 6012
rect 7728 5952 7792 5956
rect 7808 6012 7872 6016
rect 7808 5956 7812 6012
rect 7812 5956 7868 6012
rect 7868 5956 7872 6012
rect 7808 5952 7872 5956
rect 3568 5468 3632 5472
rect 3568 5412 3572 5468
rect 3572 5412 3628 5468
rect 3628 5412 3632 5468
rect 3568 5408 3632 5412
rect 3648 5468 3712 5472
rect 3648 5412 3652 5468
rect 3652 5412 3708 5468
rect 3708 5412 3712 5468
rect 3648 5408 3712 5412
rect 3728 5468 3792 5472
rect 3728 5412 3732 5468
rect 3732 5412 3788 5468
rect 3788 5412 3792 5468
rect 3728 5408 3792 5412
rect 3808 5468 3872 5472
rect 3808 5412 3812 5468
rect 3812 5412 3868 5468
rect 3868 5412 3872 5468
rect 3808 5408 3872 5412
rect 8568 5468 8632 5472
rect 8568 5412 8572 5468
rect 8572 5412 8628 5468
rect 8628 5412 8632 5468
rect 8568 5408 8632 5412
rect 8648 5468 8712 5472
rect 8648 5412 8652 5468
rect 8652 5412 8708 5468
rect 8708 5412 8712 5468
rect 8648 5408 8712 5412
rect 8728 5468 8792 5472
rect 8728 5412 8732 5468
rect 8732 5412 8788 5468
rect 8788 5412 8792 5468
rect 8728 5408 8792 5412
rect 8808 5468 8872 5472
rect 8808 5412 8812 5468
rect 8812 5412 8868 5468
rect 8868 5412 8872 5468
rect 8808 5408 8872 5412
rect 7568 4924 7632 4928
rect 7568 4868 7572 4924
rect 7572 4868 7628 4924
rect 7628 4868 7632 4924
rect 7568 4864 7632 4868
rect 7648 4924 7712 4928
rect 7648 4868 7652 4924
rect 7652 4868 7708 4924
rect 7708 4868 7712 4924
rect 7648 4864 7712 4868
rect 7728 4924 7792 4928
rect 7728 4868 7732 4924
rect 7732 4868 7788 4924
rect 7788 4868 7792 4924
rect 7728 4864 7792 4868
rect 7808 4924 7872 4928
rect 7808 4868 7812 4924
rect 7812 4868 7868 4924
rect 7868 4868 7872 4924
rect 7808 4864 7872 4868
rect 3568 4380 3632 4384
rect 3568 4324 3572 4380
rect 3572 4324 3628 4380
rect 3628 4324 3632 4380
rect 3568 4320 3632 4324
rect 3648 4380 3712 4384
rect 3648 4324 3652 4380
rect 3652 4324 3708 4380
rect 3708 4324 3712 4380
rect 3648 4320 3712 4324
rect 3728 4380 3792 4384
rect 3728 4324 3732 4380
rect 3732 4324 3788 4380
rect 3788 4324 3792 4380
rect 3728 4320 3792 4324
rect 3808 4380 3872 4384
rect 3808 4324 3812 4380
rect 3812 4324 3868 4380
rect 3868 4324 3872 4380
rect 3808 4320 3872 4324
rect 8568 4380 8632 4384
rect 8568 4324 8572 4380
rect 8572 4324 8628 4380
rect 8628 4324 8632 4380
rect 8568 4320 8632 4324
rect 8648 4380 8712 4384
rect 8648 4324 8652 4380
rect 8652 4324 8708 4380
rect 8708 4324 8712 4380
rect 8648 4320 8712 4324
rect 8728 4380 8792 4384
rect 8728 4324 8732 4380
rect 8732 4324 8788 4380
rect 8788 4324 8792 4380
rect 8728 4320 8792 4324
rect 8808 4380 8872 4384
rect 8808 4324 8812 4380
rect 8812 4324 8868 4380
rect 8868 4324 8872 4380
rect 8808 4320 8872 4324
rect 7568 3836 7632 3840
rect 7568 3780 7572 3836
rect 7572 3780 7628 3836
rect 7628 3780 7632 3836
rect 7568 3776 7632 3780
rect 7648 3836 7712 3840
rect 7648 3780 7652 3836
rect 7652 3780 7708 3836
rect 7708 3780 7712 3836
rect 7648 3776 7712 3780
rect 7728 3836 7792 3840
rect 7728 3780 7732 3836
rect 7732 3780 7788 3836
rect 7788 3780 7792 3836
rect 7728 3776 7792 3780
rect 7808 3836 7872 3840
rect 7808 3780 7812 3836
rect 7812 3780 7868 3836
rect 7868 3780 7872 3836
rect 7808 3776 7872 3780
rect 3568 3292 3632 3296
rect 3568 3236 3572 3292
rect 3572 3236 3628 3292
rect 3628 3236 3632 3292
rect 3568 3232 3632 3236
rect 3648 3292 3712 3296
rect 3648 3236 3652 3292
rect 3652 3236 3708 3292
rect 3708 3236 3712 3292
rect 3648 3232 3712 3236
rect 3728 3292 3792 3296
rect 3728 3236 3732 3292
rect 3732 3236 3788 3292
rect 3788 3236 3792 3292
rect 3728 3232 3792 3236
rect 3808 3292 3872 3296
rect 3808 3236 3812 3292
rect 3812 3236 3868 3292
rect 3868 3236 3872 3292
rect 3808 3232 3872 3236
rect 8568 3292 8632 3296
rect 8568 3236 8572 3292
rect 8572 3236 8628 3292
rect 8628 3236 8632 3292
rect 8568 3232 8632 3236
rect 8648 3292 8712 3296
rect 8648 3236 8652 3292
rect 8652 3236 8708 3292
rect 8708 3236 8712 3292
rect 8648 3232 8712 3236
rect 8728 3292 8792 3296
rect 8728 3236 8732 3292
rect 8732 3236 8788 3292
rect 8788 3236 8792 3292
rect 8728 3232 8792 3236
rect 8808 3292 8872 3296
rect 8808 3236 8812 3292
rect 8812 3236 8868 3292
rect 8868 3236 8872 3292
rect 8808 3232 8872 3236
rect 7568 2748 7632 2752
rect 7568 2692 7572 2748
rect 7572 2692 7628 2748
rect 7628 2692 7632 2748
rect 7568 2688 7632 2692
rect 7648 2748 7712 2752
rect 7648 2692 7652 2748
rect 7652 2692 7708 2748
rect 7708 2692 7712 2748
rect 7648 2688 7712 2692
rect 7728 2748 7792 2752
rect 7728 2692 7732 2748
rect 7732 2692 7788 2748
rect 7788 2692 7792 2748
rect 7728 2688 7792 2692
rect 7808 2748 7872 2752
rect 7808 2692 7812 2748
rect 7812 2692 7868 2748
rect 7868 2692 7872 2748
rect 7808 2688 7872 2692
rect 8340 2620 8404 2684
rect 3568 2204 3632 2208
rect 3568 2148 3572 2204
rect 3572 2148 3628 2204
rect 3628 2148 3632 2204
rect 3568 2144 3632 2148
rect 3648 2204 3712 2208
rect 3648 2148 3652 2204
rect 3652 2148 3708 2204
rect 3708 2148 3712 2204
rect 3648 2144 3712 2148
rect 3728 2204 3792 2208
rect 3728 2148 3732 2204
rect 3732 2148 3788 2204
rect 3788 2148 3792 2204
rect 3728 2144 3792 2148
rect 3808 2204 3872 2208
rect 3808 2148 3812 2204
rect 3812 2148 3868 2204
rect 3868 2148 3872 2204
rect 3808 2144 3872 2148
rect 8568 2204 8632 2208
rect 8568 2148 8572 2204
rect 8572 2148 8628 2204
rect 8628 2148 8632 2204
rect 8568 2144 8632 2148
rect 8648 2204 8712 2208
rect 8648 2148 8652 2204
rect 8652 2148 8708 2204
rect 8708 2148 8712 2204
rect 8648 2144 8712 2148
rect 8728 2204 8792 2208
rect 8728 2148 8732 2204
rect 8732 2148 8788 2204
rect 8788 2148 8792 2204
rect 8728 2144 8792 2148
rect 8808 2204 8872 2208
rect 8808 2148 8812 2204
rect 8812 2148 8868 2204
rect 8868 2148 8872 2204
rect 8808 2144 8872 2148
rect 8156 2076 8220 2140
rect 7568 1660 7632 1664
rect 7568 1604 7572 1660
rect 7572 1604 7628 1660
rect 7628 1604 7632 1660
rect 7568 1600 7632 1604
rect 7648 1660 7712 1664
rect 7648 1604 7652 1660
rect 7652 1604 7708 1660
rect 7708 1604 7712 1660
rect 7648 1600 7712 1604
rect 7728 1660 7792 1664
rect 7728 1604 7732 1660
rect 7732 1604 7788 1660
rect 7788 1604 7792 1660
rect 7728 1600 7792 1604
rect 7808 1660 7872 1664
rect 7808 1604 7812 1660
rect 7812 1604 7868 1660
rect 7868 1604 7872 1660
rect 7808 1600 7872 1604
rect 8156 1532 8220 1596
rect 3568 1116 3632 1120
rect 3568 1060 3572 1116
rect 3572 1060 3628 1116
rect 3628 1060 3632 1116
rect 3568 1056 3632 1060
rect 3648 1116 3712 1120
rect 3648 1060 3652 1116
rect 3652 1060 3708 1116
rect 3708 1060 3712 1116
rect 3648 1056 3712 1060
rect 3728 1116 3792 1120
rect 3728 1060 3732 1116
rect 3732 1060 3788 1116
rect 3788 1060 3792 1116
rect 3728 1056 3792 1060
rect 3808 1116 3872 1120
rect 3808 1060 3812 1116
rect 3812 1060 3868 1116
rect 3868 1060 3872 1116
rect 3808 1056 3872 1060
rect 8568 1116 8632 1120
rect 8568 1060 8572 1116
rect 8572 1060 8628 1116
rect 8628 1060 8632 1116
rect 8568 1056 8632 1060
rect 8648 1116 8712 1120
rect 8648 1060 8652 1116
rect 8652 1060 8708 1116
rect 8708 1060 8712 1116
rect 8648 1056 8712 1060
rect 8728 1116 8792 1120
rect 8728 1060 8732 1116
rect 8732 1060 8788 1116
rect 8788 1060 8792 1116
rect 8728 1056 8792 1060
rect 8808 1116 8872 1120
rect 8808 1060 8812 1116
rect 8812 1060 8868 1116
rect 8868 1060 8872 1116
rect 8808 1056 8872 1060
<< metal4 >>
rect 2560 15808 2880 15824
rect 2560 15744 2568 15808
rect 2632 15744 2648 15808
rect 2712 15744 2728 15808
rect 2792 15744 2808 15808
rect 2872 15744 2880 15808
rect 2560 14720 2880 15744
rect 2560 14656 2568 14720
rect 2632 14656 2648 14720
rect 2712 14656 2728 14720
rect 2792 14656 2808 14720
rect 2872 14656 2880 14720
rect 2560 13632 2880 14656
rect 2560 13568 2568 13632
rect 2632 13568 2648 13632
rect 2712 13568 2728 13632
rect 2792 13568 2808 13632
rect 2872 13568 2880 13632
rect 2560 13206 2880 13568
rect 2560 12970 2602 13206
rect 2838 12970 2880 13206
rect 2560 12544 2880 12970
rect 2560 12480 2568 12544
rect 2632 12480 2648 12544
rect 2712 12480 2728 12544
rect 2792 12480 2808 12544
rect 2872 12480 2880 12544
rect 1347 12340 1413 12341
rect 1347 12276 1348 12340
rect 1412 12276 1413 12340
rect 1347 12275 1413 12276
rect 1350 12069 1410 12275
rect 1347 12068 1413 12069
rect 1347 12004 1348 12068
rect 1412 12004 1413 12068
rect 1347 12003 1413 12004
rect 2560 11456 2880 12480
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9206 2880 9216
rect 2560 8970 2602 9206
rect 2838 8970 2880 9206
rect 2560 8192 2880 8970
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 7104 2880 8128
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5206 2880 5952
rect 2560 4970 2602 5206
rect 2838 4970 2880 5206
rect 2560 4893 2880 4970
rect 3560 15264 3880 15824
rect 3560 15200 3568 15264
rect 3632 15200 3648 15264
rect 3712 15200 3728 15264
rect 3792 15200 3808 15264
rect 3872 15200 3880 15264
rect 3560 14206 3880 15200
rect 3560 14176 3602 14206
rect 3838 14176 3880 14206
rect 3560 14112 3568 14176
rect 3872 14112 3880 14176
rect 3560 13970 3602 14112
rect 3838 13970 3880 14112
rect 3560 13088 3880 13970
rect 3560 13024 3568 13088
rect 3632 13024 3648 13088
rect 3712 13024 3728 13088
rect 3792 13024 3808 13088
rect 3872 13024 3880 13088
rect 3560 12000 3880 13024
rect 3560 11936 3568 12000
rect 3632 11936 3648 12000
rect 3712 11936 3728 12000
rect 3792 11936 3808 12000
rect 3872 11936 3880 12000
rect 3560 10912 3880 11936
rect 3560 10848 3568 10912
rect 3632 10848 3648 10912
rect 3712 10848 3728 10912
rect 3792 10848 3808 10912
rect 3872 10848 3880 10912
rect 3560 10206 3880 10848
rect 3560 9970 3602 10206
rect 3838 9970 3880 10206
rect 3560 9824 3880 9970
rect 3560 9760 3568 9824
rect 3632 9760 3648 9824
rect 3712 9760 3728 9824
rect 3792 9760 3808 9824
rect 3872 9760 3880 9824
rect 3560 8736 3880 9760
rect 3560 8672 3568 8736
rect 3632 8672 3648 8736
rect 3712 8672 3728 8736
rect 3792 8672 3808 8736
rect 3872 8672 3880 8736
rect 3560 7648 3880 8672
rect 3560 7584 3568 7648
rect 3632 7584 3648 7648
rect 3712 7584 3728 7648
rect 3792 7584 3808 7648
rect 3872 7584 3880 7648
rect 3560 6560 3880 7584
rect 3560 6496 3568 6560
rect 3632 6496 3648 6560
rect 3712 6496 3728 6560
rect 3792 6496 3808 6560
rect 3872 6496 3880 6560
rect 3560 6206 3880 6496
rect 3560 5970 3602 6206
rect 3838 5970 3880 6206
rect 3560 5472 3880 5970
rect 3560 5408 3568 5472
rect 3632 5408 3648 5472
rect 3712 5408 3728 5472
rect 3792 5408 3808 5472
rect 3872 5408 3880 5472
rect 3560 4384 3880 5408
rect 3560 4320 3568 4384
rect 3632 4320 3648 4384
rect 3712 4320 3728 4384
rect 3792 4320 3808 4384
rect 3872 4320 3880 4384
rect 1996 4206 2276 4248
rect 1996 3970 2018 4206
rect 2254 3970 2276 4206
rect 1996 3928 2276 3970
rect 3560 3296 3880 4320
rect 1256 3206 1536 3248
rect 1256 2970 1278 3206
rect 1514 2970 1536 3206
rect 1256 2928 1536 2970
rect 3560 3232 3568 3296
rect 3632 3232 3648 3296
rect 3712 3232 3728 3296
rect 3792 3232 3808 3296
rect 3872 3232 3880 3296
rect 3560 2208 3880 3232
rect 3560 2144 3568 2208
rect 3632 2206 3648 2208
rect 3712 2206 3728 2208
rect 3792 2206 3808 2208
rect 3872 2144 3880 2208
rect 3560 1970 3602 2144
rect 3838 1970 3880 2144
rect 3560 1120 3880 1970
rect 3560 1056 3568 1120
rect 3632 1056 3648 1120
rect 3712 1056 3728 1120
rect 3792 1056 3808 1120
rect 3872 1056 3880 1120
rect 3560 1040 3880 1056
rect 4560 15206 4880 15824
rect 4560 14970 4602 15206
rect 4838 14970 4880 15206
rect 4560 11206 4880 14970
rect 4560 10970 4602 11206
rect 4838 10970 4880 11206
rect 4560 7206 4880 10970
rect 4560 6970 4602 7206
rect 4838 6970 4880 7206
rect 4560 3206 4880 6970
rect 4560 2970 4602 3206
rect 4838 2970 4880 3206
rect 4560 1040 4880 2970
rect 5560 4206 5880 15824
rect 7560 15808 7880 15824
rect 7560 15744 7568 15808
rect 7632 15744 7648 15808
rect 7712 15744 7728 15808
rect 7792 15744 7808 15808
rect 7872 15744 7880 15808
rect 7560 14720 7880 15744
rect 7560 14656 7568 14720
rect 7632 14656 7648 14720
rect 7712 14656 7728 14720
rect 7792 14656 7808 14720
rect 7872 14656 7880 14720
rect 7235 13836 7301 13837
rect 7235 13772 7236 13836
rect 7300 13772 7301 13836
rect 7235 13771 7301 13772
rect 7238 9349 7298 13771
rect 7560 13632 7880 14656
rect 7560 13568 7568 13632
rect 7632 13568 7648 13632
rect 7712 13568 7728 13632
rect 7792 13568 7808 13632
rect 7872 13568 7880 13632
rect 7560 13206 7880 13568
rect 7560 12970 7602 13206
rect 7838 12970 7880 13206
rect 7560 12544 7880 12970
rect 7560 12480 7568 12544
rect 7632 12480 7648 12544
rect 7712 12480 7728 12544
rect 7792 12480 7808 12544
rect 7872 12480 7880 12544
rect 7560 11456 7880 12480
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 7560 10368 7880 11392
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7235 9348 7301 9349
rect 7235 9284 7236 9348
rect 7300 9284 7301 9348
rect 7235 9283 7301 9284
rect 5560 3970 5602 4206
rect 5838 3970 5880 4206
rect 5560 1040 5880 3970
rect 7560 9280 7880 10304
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 9206 7880 9216
rect 7560 8970 7602 9206
rect 7838 8970 7880 9206
rect 7560 8192 7880 8970
rect 8560 15264 8880 15824
rect 8560 15200 8568 15264
rect 8632 15200 8648 15264
rect 8712 15200 8728 15264
rect 8792 15200 8808 15264
rect 8872 15200 8880 15264
rect 8560 14206 8880 15200
rect 8560 14176 8602 14206
rect 8838 14176 8880 14206
rect 8560 14112 8568 14176
rect 8872 14112 8880 14176
rect 8560 13970 8602 14112
rect 8838 13970 8880 14112
rect 8560 13088 8880 13970
rect 8560 13024 8568 13088
rect 8632 13024 8648 13088
rect 8712 13024 8728 13088
rect 8792 13024 8808 13088
rect 8872 13024 8880 13088
rect 8560 12000 8880 13024
rect 8560 11936 8568 12000
rect 8632 11936 8648 12000
rect 8712 11936 8728 12000
rect 8792 11936 8808 12000
rect 8872 11936 8880 12000
rect 8560 10912 8880 11936
rect 8560 10848 8568 10912
rect 8632 10848 8648 10912
rect 8712 10848 8728 10912
rect 8792 10848 8808 10912
rect 8872 10848 8880 10912
rect 8560 10206 8880 10848
rect 8560 9970 8602 10206
rect 8838 9970 8880 10206
rect 8560 9824 8880 9970
rect 8560 9760 8568 9824
rect 8632 9760 8648 9824
rect 8712 9760 8728 9824
rect 8792 9760 8808 9824
rect 8872 9760 8880 9824
rect 8339 8940 8405 8941
rect 8339 8876 8340 8940
rect 8404 8876 8405 8940
rect 8339 8875 8405 8876
rect 7560 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7880 8192
rect 7560 7104 7880 8128
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 6016 7880 7040
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 5206 7880 5952
rect 7560 4970 7602 5206
rect 7838 4970 7880 5206
rect 7560 4928 7880 4970
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 7560 3840 7880 4864
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 2752 7880 3776
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 1664 7880 2688
rect 8342 2685 8402 8875
rect 8560 8736 8880 9760
rect 8560 8672 8568 8736
rect 8632 8672 8648 8736
rect 8712 8672 8728 8736
rect 8792 8672 8808 8736
rect 8872 8672 8880 8736
rect 8560 7648 8880 8672
rect 8560 7584 8568 7648
rect 8632 7584 8648 7648
rect 8712 7584 8728 7648
rect 8792 7584 8808 7648
rect 8872 7584 8880 7648
rect 8560 6560 8880 7584
rect 8560 6496 8568 6560
rect 8632 6496 8648 6560
rect 8712 6496 8728 6560
rect 8792 6496 8808 6560
rect 8872 6496 8880 6560
rect 8560 6206 8880 6496
rect 8560 5970 8602 6206
rect 8838 5970 8880 6206
rect 8560 5472 8880 5970
rect 8560 5408 8568 5472
rect 8632 5408 8648 5472
rect 8712 5408 8728 5472
rect 8792 5408 8808 5472
rect 8872 5408 8880 5472
rect 8560 4384 8880 5408
rect 8560 4320 8568 4384
rect 8632 4320 8648 4384
rect 8712 4320 8728 4384
rect 8792 4320 8808 4384
rect 8872 4320 8880 4384
rect 8560 3296 8880 4320
rect 8560 3232 8568 3296
rect 8632 3232 8648 3296
rect 8712 3232 8728 3296
rect 8792 3232 8808 3296
rect 8872 3232 8880 3296
rect 8339 2684 8405 2685
rect 8339 2620 8340 2684
rect 8404 2620 8405 2684
rect 8339 2619 8405 2620
rect 8560 2208 8880 3232
rect 8560 2144 8568 2208
rect 8632 2206 8648 2208
rect 8712 2206 8728 2208
rect 8792 2206 8808 2208
rect 8872 2144 8880 2208
rect 8155 2140 8221 2141
rect 8155 2076 8156 2140
rect 8220 2076 8221 2140
rect 8155 2075 8221 2076
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 7560 1206 7880 1600
rect 8158 1597 8218 2075
rect 8560 1970 8602 2144
rect 8838 1970 8880 2144
rect 8155 1596 8221 1597
rect 8155 1532 8156 1596
rect 8220 1532 8221 1596
rect 8155 1531 8221 1532
rect 7560 970 7602 1206
rect 7838 970 7880 1206
rect 8560 1120 8880 1970
rect 8560 1056 8568 1120
rect 8632 1056 8648 1120
rect 8712 1056 8728 1120
rect 8792 1056 8808 1120
rect 8872 1056 8880 1120
rect 8560 1040 8880 1056
rect 9560 15206 9880 15824
rect 9560 14970 9602 15206
rect 9838 14970 9880 15206
rect 9560 11206 9880 14970
rect 9560 10970 9602 11206
rect 9838 10970 9880 11206
rect 9560 7206 9880 10970
rect 9560 6970 9602 7206
rect 9838 6970 9880 7206
rect 9560 3206 9880 6970
rect 9560 2970 9602 3206
rect 9838 2970 9880 3206
rect 9560 1040 9880 2970
rect 7560 928 7880 970
<< via4 >>
rect 2602 12970 2838 13206
rect 2602 8970 2838 9206
rect 2602 4970 2838 5206
rect 3602 14176 3838 14206
rect 3602 14112 3632 14176
rect 3632 14112 3648 14176
rect 3648 14112 3712 14176
rect 3712 14112 3728 14176
rect 3728 14112 3792 14176
rect 3792 14112 3808 14176
rect 3808 14112 3838 14176
rect 3602 13970 3838 14112
rect 3602 9970 3838 10206
rect 3602 5970 3838 6206
rect 2018 3970 2254 4206
rect 1278 2970 1514 3206
rect 3602 2144 3632 2206
rect 3632 2144 3648 2206
rect 3648 2144 3712 2206
rect 3712 2144 3728 2206
rect 3728 2144 3792 2206
rect 3792 2144 3808 2206
rect 3808 2144 3838 2206
rect 3602 1970 3838 2144
rect 4602 14970 4838 15206
rect 4602 10970 4838 11206
rect 4602 6970 4838 7206
rect 4602 2970 4838 3206
rect 7602 12970 7838 13206
rect 5602 3970 5838 4206
rect 7602 8970 7838 9206
rect 8602 14176 8838 14206
rect 8602 14112 8632 14176
rect 8632 14112 8648 14176
rect 8648 14112 8712 14176
rect 8712 14112 8728 14176
rect 8728 14112 8792 14176
rect 8792 14112 8808 14176
rect 8808 14112 8838 14176
rect 8602 13970 8838 14112
rect 8602 9970 8838 10206
rect 7602 4970 7838 5206
rect 8602 5970 8838 6206
rect 8602 2144 8632 2206
rect 8632 2144 8648 2206
rect 8648 2144 8712 2206
rect 8712 2144 8728 2206
rect 8728 2144 8792 2206
rect 8792 2144 8808 2206
rect 8808 2144 8838 2206
rect 8602 1970 8838 2144
rect 7602 970 7838 1206
rect 9602 14970 9838 15206
rect 9602 10970 9838 11206
rect 9602 6970 9838 7206
rect 9602 2970 9838 3206
<< metal5 >>
rect 872 15206 9892 15248
rect 872 14970 4602 15206
rect 4838 14970 9602 15206
rect 9838 14970 9892 15206
rect 872 14928 9892 14970
rect 872 14206 9892 14248
rect 872 13970 3602 14206
rect 3838 13970 8602 14206
rect 8838 13970 9892 14206
rect 872 13928 9892 13970
rect 872 13206 9892 13248
rect 872 12970 2602 13206
rect 2838 12970 7602 13206
rect 7838 12970 9892 13206
rect 872 12928 9892 12970
rect 872 11206 9892 11248
rect 872 10970 4602 11206
rect 4838 10970 9602 11206
rect 9838 10970 9892 11206
rect 872 10928 9892 10970
rect 872 10206 9892 10248
rect 872 9970 3602 10206
rect 3838 9970 8602 10206
rect 8838 9970 9892 10206
rect 872 9928 9892 9970
rect 872 9206 9892 9248
rect 872 8970 2602 9206
rect 2838 8970 7602 9206
rect 7838 8970 9892 9206
rect 872 8928 9892 8970
rect 872 7206 9892 7248
rect 872 6970 4602 7206
rect 4838 6970 9602 7206
rect 9838 6970 9892 7206
rect 872 6928 9892 6970
rect 872 6206 9892 6248
rect 872 5970 3602 6206
rect 3838 5970 8602 6206
rect 8838 5970 9892 6206
rect 872 5928 9892 5970
rect 872 5206 9892 5248
rect 872 4970 2602 5206
rect 2838 4970 7602 5206
rect 7838 4970 9892 5206
rect 872 4928 9892 4970
rect 872 4206 9892 4248
rect 872 3970 2018 4206
rect 2254 3970 5602 4206
rect 5838 3970 9892 4206
rect 872 3928 9892 3970
rect 872 3206 9892 3248
rect 872 2970 1278 3206
rect 1514 2970 4602 3206
rect 4838 2970 9602 3206
rect 9838 2970 9892 3206
rect 872 2928 9892 2970
rect 872 2206 9892 2248
rect 872 1970 3602 2206
rect 3838 1970 8602 2206
rect 8838 1970 9892 2206
rect 872 1928 9892 1970
rect 872 1206 9892 1248
rect 872 970 7602 1206
rect 7838 970 9892 1206
rect 872 928 9892 970
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 3312 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 3772 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1663720911
transform 1 0 4416 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 5060 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52
timestamp 1663720911
transform 1 0 5704 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1663720911
transform 1 0 6164 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64
timestamp 1663720911
transform 1 0 6808 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 7452 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 8280 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92
timestamp 1663720911
transform 1 0 9384 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1663720911
transform 1 0 3312 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_31
timestamp 1663720911
transform 1 0 3772 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1663720911
transform 1 0 4416 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1663720911
transform 1 0 5060 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1663720911
transform 1 0 5704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_59
timestamp 1663720911
transform 1 0 6348 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_66
timestamp 1663720911
transform 1 0 6992 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_73
timestamp 1663720911
transform 1 0 7636 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_80
timestamp 1663720911
transform 1 0 8280 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 1663720911
transform 1 0 8740 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1663720911
transform 1 0 9384 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1663720911
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_31
timestamp 1663720911
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 1663720911
transform 1 0 4508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_44
timestamp 1663720911
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 5520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_52
timestamp 1663720911
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1663720911
transform 1 0 6164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 1663720911
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_71
timestamp 1663720911
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_79 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1663720911
transform 1 0 8740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_92
timestamp 1663720911
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1663720911
transform 1 0 3312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1663720911
transform 1 0 4324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_44
timestamp 1663720911
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1663720911
transform 1 0 5612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_58
timestamp 1663720911
transform 1 0 6256 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1663720911
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_76
timestamp 1663720911
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_80
timestamp 1663720911
transform 1 0 8280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1663720911
transform 1 0 8740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1663720911
transform 1 0 9384 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1663720911
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_31
timestamp 1663720911
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_38
timestamp 1663720911
transform 1 0 4416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_42
timestamp 1663720911
transform 1 0 4784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_46
timestamp 1663720911
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_50
timestamp 1663720911
transform 1 0 5520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_52
timestamp 1663720911
transform 1 0 5704 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_57
timestamp 1663720911
transform 1 0 6164 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_65
timestamp 1663720911
transform 1 0 6900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_69
timestamp 1663720911
transform 1 0 7268 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 1663720911
transform 1 0 8004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_82
timestamp 1663720911
transform 1 0 8464 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_92
timestamp 1663720911
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_26
timestamp 1663720911
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1663720911
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1663720911
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1663720911
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_59
timestamp 1663720911
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp 1663720911
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_67
timestamp 1663720911
transform 1 0 7084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_74
timestamp 1663720911
transform 1 0 7728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_78
timestamp 1663720911
transform 1 0 8096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_80
timestamp 1663720911
transform 1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1663720911
transform 1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1663720911
transform 1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_31
timestamp 1663720911
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 1663720911
transform 1 0 4784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_49
timestamp 1663720911
transform 1 0 5428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_52
timestamp 1663720911
transform 1 0 5704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1663720911
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_65
timestamp 1663720911
transform 1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_72
timestamp 1663720911
transform 1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp 1663720911
transform 1 0 8280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_84
timestamp 1663720911
transform 1 0 8648 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_92
timestamp 1663720911
transform 1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_26
timestamp 1663720911
transform 1 0 3312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_32
timestamp 1663720911
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_36
timestamp 1663720911
transform 1 0 4232 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_44
timestamp 1663720911
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_54
timestamp 1663720911
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_58
timestamp 1663720911
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_64
timestamp 1663720911
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_71
timestamp 1663720911
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_80
timestamp 1663720911
transform 1 0 8280 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_86
timestamp 1663720911
transform 1 0 8832 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_91
timestamp 1663720911
transform 1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1663720911
transform 1 0 1196 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_10
timestamp 1663720911
transform 1 0 1840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_18
timestamp 1663720911
transform 1 0 2576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1663720911
transform 1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1663720911
transform 1 0 3588 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1663720911
transform 1 0 5612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_55
timestamp 1663720911
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_57
timestamp 1663720911
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_67
timestamp 1663720911
transform 1 0 7084 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_75
timestamp 1663720911
transform 1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1663720911
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1663720911
transform 1 0 8740 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_91
timestamp 1663720911
transform 1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1663720911
transform 1 0 1196 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1663720911
transform 1 0 1564 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_16
timestamp 1663720911
transform 1 0 2392 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_24
timestamp 1663720911
transform 1 0 3128 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1663720911
transform 1 0 5060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_49
timestamp 1663720911
transform 1 0 5428 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1663720911
transform 1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1663720911
transform 1 0 6164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_87
timestamp 1663720911
transform 1 0 8924 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_93
timestamp 1663720911
transform 1 0 9476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1663720911
transform 1 0 1196 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1663720911
transform 1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1663720911
transform 1 0 3588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_52
timestamp 1663720911
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1663720911
transform 1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1663720911
transform 1 0 8740 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_92
timestamp 1663720911
transform 1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1663720911
transform 1 0 1196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1663720911
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1663720911
transform 1 0 3680 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1663720911
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1663720911
transform 1 0 6164 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1663720911
transform 1 0 8740 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1663720911
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1663720911
transform 1 0 1196 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1663720911
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1663720911
transform 1 0 3588 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_39
timestamp 1663720911
transform 1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_67
timestamp 1663720911
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1663720911
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1663720911
transform 1 0 8556 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1663720911
transform 1 0 8740 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_92
timestamp 1663720911
transform 1 0 9384 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1663720911
transform 1 0 1196 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1663720911
transform 1 0 1564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_16
timestamp 1663720911
transform 1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_46
timestamp 1663720911
transform 1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1663720911
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1663720911
transform 1 0 6164 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_67
timestamp 1663720911
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp 1663720911
transform 1 0 9384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1663720911
transform 1 0 1196 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1663720911
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1663720911
transform 1 0 3588 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp 1663720911
transform 1 0 3956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_42
timestamp 1663720911
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1663720911
transform 1 0 5152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_67
timestamp 1663720911
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1663720911
transform 1 0 8004 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1663720911
transform 1 0 8556 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1663720911
transform 1 0 8740 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_91
timestamp 1663720911
transform 1 0 9292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1663720911
transform 1 0 1196 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1663720911
transform 1 0 3128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1663720911
transform 1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1663720911
transform 1 0 6164 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 1663720911
transform 1 0 6992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_90
timestamp 1663720911
transform 1 0 9200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1663720911
transform 1 0 1196 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_14
timestamp 1663720911
transform 1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1663720911
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1663720911
transform 1 0 3588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_51
timestamp 1663720911
transform 1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1663720911
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1663720911
transform 1 0 8740 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_92
timestamp 1663720911
transform 1 0 9384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1663720911
transform 1 0 1196 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1663720911
transform 1 0 2116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_43
timestamp 1663720911
transform 1 0 4876 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1663720911
transform 1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1663720911
transform 1 0 6164 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1663720911
transform 1 0 8740 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_92
timestamp 1663720911
transform 1 0 9384 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1663720911
transform 1 0 1196 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1663720911
transform 1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1663720911
transform 1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1663720911
transform 1 0 3588 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_45
timestamp 1663720911
transform 1 0 5060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 1663720911
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1663720911
transform 1 0 8096 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1663720911
transform 1 0 8740 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_91
timestamp 1663720911
transform 1 0 9292 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1663720911
transform 1 0 1196 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 1663720911
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_30
timestamp 1663720911
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1663720911
transform 1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1663720911
transform 1 0 6164 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_79
timestamp 1663720911
transform 1 0 8188 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_91
timestamp 1663720911
transform 1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1663720911
transform 1 0 1196 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1663720911
transform 1 0 3312 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1663720911
transform 1 0 3588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 1663720911
transform 1 0 4048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_64
timestamp 1663720911
transform 1 0 6808 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_70
timestamp 1663720911
transform 1 0 7360 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1663720911
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1663720911
transform 1 0 8556 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1663720911
transform 1 0 8740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_92
timestamp 1663720911
transform 1 0 9384 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1663720911
transform 1 0 1196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_14
timestamp 1663720911
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_44
timestamp 1663720911
transform 1 0 4968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1663720911
transform 1 0 5888 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1663720911
transform 1 0 6164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_81
timestamp 1663720911
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_85
timestamp 1663720911
transform 1 0 8740 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp 1663720911
transform 1 0 9384 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1663720911
transform 1 0 1196 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1663720911
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1663720911
transform 1 0 3588 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_40
timestamp 1663720911
transform 1 0 4600 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_72
timestamp 1663720911
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_76
timestamp 1663720911
transform 1 0 7912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1663720911
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1663720911
transform 1 0 8740 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_91
timestamp 1663720911
transform 1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1663720911
transform 1 0 1196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_14
timestamp 1663720911
transform 1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_44
timestamp 1663720911
transform 1 0 4968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_48
timestamp 1663720911
transform 1 0 5336 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1663720911
transform 1 0 5888 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1663720911
transform 1 0 6164 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1663720911
transform 1 0 6532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_88
timestamp 1663720911
transform 1 0 9016 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1663720911
transform 1 0 1196 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1663720911
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1663720911
transform 1 0 3588 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_34
timestamp 1663720911
transform 1 0 4048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_43
timestamp 1663720911
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_67
timestamp 1663720911
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1663720911
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1663720911
transform 1 0 8740 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_92
timestamp 1663720911
transform 1 0 9384 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1663720911
transform 1 0 1196 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_11
timestamp 1663720911
transform 1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1663720911
transform 1 0 2300 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1663720911
transform 1 0 2852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 1663720911
transform 1 0 3680 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_42
timestamp 1663720911
transform 1 0 4784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1663720911
transform 1 0 5888 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1663720911
transform 1 0 6164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_61
timestamp 1663720911
transform 1 0 6532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_82
timestamp 1663720911
transform 1 0 8464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_86
timestamp 1663720911
transform 1 0 8832 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_91
timestamp 1663720911
transform 1 0 9292 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1663720911
transform 1 0 1196 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_10
timestamp 1663720911
transform 1 0 1840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_18
timestamp 1663720911
transform 1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1663720911
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1663720911
transform 1 0 3588 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_46
timestamp 1663720911
transform 1 0 5152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_54
timestamp 1663720911
transform 1 0 5888 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_57
timestamp 1663720911
transform 1 0 6164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 1663720911
transform 1 0 6532 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1663720911
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1663720911
transform 1 0 8740 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_91
timestamp 1663720911
transform 1 0 9292 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1663720911
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1663720911
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1663720911
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1663720911
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1663720911
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1663720911
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1663720911
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1663720911
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1663720911
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1663720911
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1663720911
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1663720911
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1663720911
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1663720911
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1663720911
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1663720911
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1663720911
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1663720911
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1663720911
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1663720911
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1663720911
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1663720911
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1663720911
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1663720911
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1663720911
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1663720911
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1663720911
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1663720911
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1663720911
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1663720911
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1663720911
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1663720911
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1663720911
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1663720911
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1663720911
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1663720911
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1663720911
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1663720911
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1663720911
transform 1 0 920 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1663720911
transform -1 0 9844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1663720911
transform 1 0 920 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1663720911
transform -1 0 9844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1663720911
transform 1 0 920 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1663720911
transform -1 0 9844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1663720911
transform 1 0 920 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1663720911
transform -1 0 9844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1663720911
transform 1 0 920 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1663720911
transform -1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1663720911
transform 1 0 920 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1663720911
transform -1 0 9844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1663720911
transform 1 0 920 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1663720911
transform -1 0 9844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1663720911
transform 1 0 920 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1663720911
transform -1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1663720911
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1663720911
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1663720911
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1663720911
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1663720911
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1663720911
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1663720911
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1663720911
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1663720911
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1663720911
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1663720911
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1663720911
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1663720911
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1663720911
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1663720911
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1663720911
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1663720911
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1663720911
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1663720911
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1663720911
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1663720911
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1663720911
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1663720911
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1663720911
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1663720911
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1663720911
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1663720911
transform 1 0 6072 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1663720911
transform 1 0 3496 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1663720911
transform 1 0 8648 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1663720911
transform 1 0 6072 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1663720911
transform 1 0 3496 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1663720911
transform 1 0 8648 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1663720911
transform 1 0 6072 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1663720911
transform 1 0 3496 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1663720911
transform 1 0 8648 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1663720911
transform 1 0 6072 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1663720911
transform 1 0 3496 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1663720911
transform 1 0 6072 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1663720911
transform 1 0 8648 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 6440 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 6808 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 9384 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 9292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _090_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1663720911
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _093_
timestamp 1663720911
transform -1 0 6992 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 8924 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1663720911
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _097_
timestamp 1663720911
transform -1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _098_
timestamp 1663720911
transform 1 0 2944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _099_
timestamp 1663720911
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _100_
timestamp 1663720911
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1663720911
transform -1 0 9384 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 2392 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 5336 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _106__5
timestamp 1663720911
transform -1 0 6164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp 1663720911
transform -1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _108_
timestamp 1663720911
transform 1 0 7452 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _109_
timestamp 1663720911
transform 1 0 4784 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _110_
timestamp 1663720911
transform 1 0 1472 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1663720911
transform -1 0 4416 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112__6
timestamp 1663720911
transform -1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _113_
timestamp 1663720911
transform 1 0 6072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _114_
timestamp 1663720911
transform -1 0 4876 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1663720911
transform -1 0 4784 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116__7
timestamp 1663720911
transform 1 0 3496 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _117_
timestamp 1663720911
transform -1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _118_
timestamp 1663720911
transform -1 0 5888 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1663720911
transform -1 0 5704 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120__8
timestamp 1663720911
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _121_
timestamp 1663720911
transform 1 0 6072 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 1663720911
transform 1 0 7636 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1663720911
transform -1 0 3772 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124__9
timestamp 1663720911
transform -1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _125_
timestamp 1663720911
transform 1 0 5888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _126_
timestamp 1663720911
transform 1 0 1380 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1663720911
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _128__10
timestamp 1663720911
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _129_
timestamp 1663720911
transform 1 0 3496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _130_
timestamp 1663720911
transform 1 0 3220 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1663720911
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _132__11
timestamp 1663720911
transform 1 0 7360 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _133_
timestamp 1663720911
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _134_
timestamp 1663720911
transform 1 0 5428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1663720911
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136__12
timestamp 1663720911
transform -1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _137_
timestamp 1663720911
transform -1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _138_
timestamp 1663720911
transform 1 0 8924 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1663720911
transform -1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _140__13
timestamp 1663720911
transform 1 0 9108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _141_
timestamp 1663720911
transform 1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _142_
timestamp 1663720911
transform 1 0 8924 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1663720911
transform -1 0 6256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144__14
timestamp 1663720911
transform 1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _145_
timestamp 1663720911
transform 1 0 6992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _146_
timestamp 1663720911
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1663720911
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148__1
timestamp 1663720911
transform -1 0 4232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _149_
timestamp 1663720911
transform 1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _150_
timestamp 1663720911
transform 1 0 8924 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1663720911
transform -1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _152__2
timestamp 1663720911
transform -1 0 6900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _153_
timestamp 1663720911
transform 1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _154_
timestamp 1663720911
transform 1 0 8924 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1663720911
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156__3
timestamp 1663720911
transform 1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _157_
timestamp 1663720911
transform 1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _158__4
timestamp 1663720911
transform 1 0 4784 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 4968 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _160_
timestamp 1663720911
transform 1 0 2484 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _161_
timestamp 1663720911
transform 1 0 4416 0 1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _162_
timestamp 1663720911
transform 1 0 5152 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _163_
timestamp 1663720911
transform 1 0 2760 0 -1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _164_
timestamp 1663720911
transform 1 0 3496 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _165_
timestamp 1663720911
transform 1 0 2576 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _166_
timestamp 1663720911
transform 1 0 5980 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _167_
timestamp 1663720911
transform -1 0 8740 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _168_
timestamp 1663720911
transform -1 0 9016 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _169_
timestamp 1663720911
transform 1 0 6348 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _170_
timestamp 1663720911
transform 1 0 6072 0 1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _171_
timestamp 1663720911
transform 1 0 6532 0 -1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__dfrtp_1  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 8464 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _173_
timestamp 1663720911
transform -1 0 3312 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _174_
timestamp 1663720911
transform -1 0 3312 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _175_
timestamp 1663720911
transform 1 0 1472 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _176_
timestamp 1663720911
transform 1 0 1472 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _177_
timestamp 1663720911
transform 1 0 3772 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _178_
timestamp 1663720911
transform -1 0 5704 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _179_
timestamp 1663720911
transform 1 0 4048 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _180_
timestamp 1663720911
transform -1 0 5060 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _181_
timestamp 1663720911
transform -1 0 3680 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _182_
timestamp 1663720911
transform 1 0 3772 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _183_
timestamp 1663720911
transform 1 0 6348 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _184_
timestamp 1663720911
transform 1 0 6532 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _185_
timestamp 1663720911
transform -1 0 8464 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 1663720911
transform -1 0 4416 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 2576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _188_
timestamp 1663720911
transform -1 0 1840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_8  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 9384 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 5888 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock
timestamp 1663720911
transform -1 0 7268 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 1663720911
transform -1 0 9200 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__068_
timestamp 1663720911
transform 1 0 1472 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_clock
timestamp 1663720911
transform -1 0 3680 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_load
timestamp 1663720911
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__068_
timestamp 1663720911
transform 1 0 1472 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_clock
timestamp 1663720911
transform 1 0 5244 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_load
timestamp 1663720911
transform -1 0 7084 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 8740 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1663720911
transform -1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 9384 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 1472 0 -1 9792
box -38 -48 1694 592
use gpio_logic_high  gpio_logic_high
timestamp 0
transform 1 0 1196 0 1 1680
box -1196 -1680 32804 15320
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1663720911
transform 1 0 1472 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1663720911
transform 1 0 1656 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1663720911
transform 1 0 4048 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1663720911
transform 1 0 1656 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1663720911
transform 1 0 7636 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1663720911
transform 1 0 7452 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1663720911
transform 1 0 1472 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1663720911
transform 1 0 4048 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1663720911
transform 1 0 1472 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1663720911
transform 1 0 6348 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1663720911
transform 1 0 5152 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1663720911
transform -1 0 8188 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1663720911
transform -1 0 5888 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1663720911
transform 1 0 1472 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1663720911
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1663720911
transform 1 0 2576 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1663720911
transform 1 0 2576 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1663720911
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1663720911
transform 1 0 4324 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output1
timestamp 1663720911
transform 1 0 9016 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 1663720911
transform -1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1663720911
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1663720911
transform 1 0 9016 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1663720911
transform -1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1663720911
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1663720911
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1663720911
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1663720911
transform -1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1663720911
transform 1 0 8924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1663720911
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1663720911
transform -1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1663720911
transform 1 0 8004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1663720911
transform 1 0 5520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  output15
timestamp 1663720911
transform 1 0 3588 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output16
timestamp 1663720911
transform -1 0 5152 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output17
timestamp 1663720911
transform 1 0 3496 0 -1 3264
box -38 -48 866 592
<< labels >>
flabel metal2 s 938 16200 994 17000 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 0 nsew signal input
flabel metal2 s 5538 16200 5594 17000 0 FreeSans 224 90 0 0 gpio_defaults[10]
port 1 nsew signal input
flabel metal2 s 5998 16200 6054 17000 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 2 nsew signal input
flabel metal2 s 6458 16200 6514 17000 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 3 nsew signal input
flabel metal2 s 1398 16200 1454 17000 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 4 nsew signal input
flabel metal2 s 1858 16200 1914 17000 0 FreeSans 224 90 0 0 gpio_defaults[2]
port 5 nsew signal input
flabel metal2 s 2318 16200 2374 17000 0 FreeSans 224 90 0 0 gpio_defaults[3]
port 6 nsew signal input
flabel metal2 s 2778 16200 2834 17000 0 FreeSans 224 90 0 0 gpio_defaults[4]
port 7 nsew signal input
flabel metal2 s 3238 16200 3294 17000 0 FreeSans 224 90 0 0 gpio_defaults[5]
port 8 nsew signal input
flabel metal2 s 3698 16200 3754 17000 0 FreeSans 224 90 0 0 gpio_defaults[6]
port 9 nsew signal input
flabel metal2 s 4158 16200 4214 17000 0 FreeSans 224 90 0 0 gpio_defaults[7]
port 10 nsew signal input
flabel metal2 s 4618 16200 4674 17000 0 FreeSans 224 90 0 0 gpio_defaults[8]
port 11 nsew signal input
flabel metal2 s 5078 16200 5134 17000 0 FreeSans 224 90 0 0 gpio_defaults[9]
port 12 nsew signal input
flabel metal3 s 14000 4904 34000 5024 0 FreeSans 480 0 0 0 mgmt_gpio_in
port 13 nsew signal tristate
flabel metal3 s 14000 5720 34000 5840 0 FreeSans 480 0 0 0 mgmt_gpio_oeb
port 14 nsew signal input
flabel metal3 s 14000 6128 34000 6248 0 FreeSans 480 0 0 0 mgmt_gpio_out
port 15 nsew signal input
flabel metal3 s 14000 5312 34000 5432 0 FreeSans 480 0 0 0 one
port 16 nsew signal tristate
flabel metal3 s 14000 6536 34000 6656 0 FreeSans 480 0 0 0 pad_gpio_ana_en
port 17 nsew signal tristate
flabel metal3 s 14000 6944 34000 7064 0 FreeSans 480 0 0 0 pad_gpio_ana_pol
port 18 nsew signal tristate
flabel metal3 s 14000 7352 34000 7472 0 FreeSans 480 0 0 0 pad_gpio_ana_sel
port 19 nsew signal tristate
flabel metal3 s 14000 7760 34000 7880 0 FreeSans 480 0 0 0 pad_gpio_dm[0]
port 20 nsew signal tristate
flabel metal3 s 14000 8168 34000 8288 0 FreeSans 480 0 0 0 pad_gpio_dm[1]
port 21 nsew signal tristate
flabel metal3 s 14000 8576 34000 8696 0 FreeSans 480 0 0 0 pad_gpio_dm[2]
port 22 nsew signal tristate
flabel metal3 s 14000 8984 34000 9104 0 FreeSans 480 0 0 0 pad_gpio_holdover
port 23 nsew signal tristate
flabel metal3 s 14000 9392 34000 9512 0 FreeSans 480 0 0 0 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
flabel metal3 s 14000 9800 34000 9920 0 FreeSans 480 0 0 0 pad_gpio_in
port 25 nsew signal input
flabel metal3 s 14000 10208 34000 10328 0 FreeSans 480 0 0 0 pad_gpio_inenb
port 26 nsew signal tristate
flabel metal3 s 14000 10616 34000 10736 0 FreeSans 480 0 0 0 pad_gpio_out
port 27 nsew signal tristate
flabel metal3 s 14000 11024 34000 11144 0 FreeSans 480 0 0 0 pad_gpio_outenb
port 28 nsew signal tristate
flabel metal3 s 14000 11432 34000 11552 0 FreeSans 480 0 0 0 pad_gpio_slow_sel
port 29 nsew signal tristate
flabel metal3 s 14000 11840 34000 11960 0 FreeSans 480 0 0 0 pad_gpio_vtrip_sel
port 30 nsew signal tristate
flabel metal3 s 14000 12248 34000 12368 0 FreeSans 480 0 0 0 resetn
port 31 nsew signal input
flabel metal3 s 14000 12656 34000 12776 0 FreeSans 480 0 0 0 resetn_out
port 32 nsew signal tristate
flabel metal3 s 14000 13064 34000 13184 0 FreeSans 480 0 0 0 serial_clock
port 33 nsew signal input
flabel metal3 s 14000 13472 34000 13592 0 FreeSans 480 0 0 0 serial_clock_out
port 34 nsew signal tristate
flabel metal3 s 14000 13880 34000 14000 0 FreeSans 480 0 0 0 serial_data_in
port 35 nsew signal input
flabel metal3 s 14000 14288 34000 14408 0 FreeSans 480 0 0 0 serial_data_out
port 36 nsew signal tristate
flabel metal3 s 14000 14696 34000 14816 0 FreeSans 480 0 0 0 serial_load
port 37 nsew signal input
flabel metal3 s 14000 15104 34000 15224 0 FreeSans 480 0 0 0 serial_load_out
port 38 nsew signal tristate
flabel metal3 s 14000 15512 34000 15632 0 FreeSans 480 0 0 0 user_gpio_in
port 39 nsew signal tristate
flabel metal3 s 14000 15920 34000 16040 0 FreeSans 480 0 0 0 user_gpio_oeb
port 40 nsew signal input
flabel metal3 s 14000 16328 34000 16448 0 FreeSans 480 0 0 0 user_gpio_out
port 41 nsew signal input
flabel metal4 s 2560 4893 2880 15824 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 7560 928 7880 15824 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 928 9892 1248 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 4928 9892 5248 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 8928 9892 9248 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 12928 9892 13248 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 4560 1040 4880 15824 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 9560 1040 9880 15824 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 2928 9892 3248 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 6928 9892 7248 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 10928 9892 11248 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 14928 9892 15248 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 3560 1040 3880 15824 0 FreeSans 1920 90 0 0 vssd
port 44 nsew ground bidirectional
flabel metal4 s 8560 1040 8880 15824 0 FreeSans 1920 90 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 1928 9892 2248 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 5928 9892 6248 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 9928 9892 10248 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 13928 9892 14248 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal4 s 5560 1040 5880 15824 0 FreeSans 1920 90 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 3928 9892 4248 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal3 s 14000 4496 34000 4616 0 FreeSans 480 0 0 0 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 17000
<< end >>
