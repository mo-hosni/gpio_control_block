magic
tech sky130A
magscale 1 2
timestamp 1664316535
<< viali >>
rect 3249 15657 3283 15691
rect 9137 15657 9171 15691
rect 5457 15521 5491 15555
rect 8125 15521 8159 15555
rect 1777 15453 1811 15487
rect 4077 15453 4111 15487
rect 5733 15453 5767 15487
rect 8401 15453 8435 15487
rect 8953 15453 8987 15487
rect 2881 15385 2915 15419
rect 3065 15385 3099 15419
rect 4629 15385 4663 15419
rect 1593 15317 1627 15351
rect 6653 15317 6687 15351
rect 6653 15113 6687 15147
rect 2053 15045 2087 15079
rect 3249 15045 3283 15079
rect 8125 15045 8159 15079
rect 1409 14977 1443 15011
rect 2237 14977 2271 15011
rect 3065 14977 3099 15011
rect 9045 14977 9079 15011
rect 3801 14909 3835 14943
rect 4353 14909 4387 14943
rect 5365 14909 5399 14943
rect 8401 14909 8435 14943
rect 2421 14841 2455 14875
rect 4813 14841 4847 14875
rect 1501 14773 1535 14807
rect 2881 14773 2915 14807
rect 9229 14773 9263 14807
rect 4169 14569 4203 14603
rect 3249 14433 3283 14467
rect 4813 14433 4847 14467
rect 8125 14365 8159 14399
rect 2973 14297 3007 14331
rect 7021 14297 7055 14331
rect 8953 14297 8987 14331
rect 9137 14297 9171 14331
rect 1501 14229 1535 14263
rect 5549 14229 5583 14263
rect 7481 14229 7515 14263
rect 9321 14229 9355 14263
rect 5733 14025 5767 14059
rect 5549 13957 5583 13991
rect 2605 13889 2639 13923
rect 4445 13889 4479 13923
rect 5365 13889 5399 13923
rect 6653 13889 6687 13923
rect 7021 13889 7055 13923
rect 8493 13889 8527 13923
rect 1593 13821 1627 13855
rect 2145 13821 2179 13855
rect 2973 13821 3007 13855
rect 4905 13821 4939 13855
rect 8953 13821 8987 13855
rect 7481 13481 7515 13515
rect 4445 13345 4479 13379
rect 5549 13345 5583 13379
rect 3893 13277 3927 13311
rect 5181 13277 5215 13311
rect 7021 13277 7055 13311
rect 8033 13277 8067 13311
rect 8953 13277 8987 13311
rect 1501 13209 1535 13243
rect 2789 13141 2823 13175
rect 8217 13141 8251 13175
rect 9137 13141 9171 13175
rect 8309 12937 8343 12971
rect 1501 12801 1535 12835
rect 2881 12801 2915 12835
rect 4353 12801 4387 12835
rect 5365 12801 5399 12835
rect 9229 12801 9263 12835
rect 2513 12733 2547 12767
rect 5641 12733 5675 12767
rect 6561 12733 6595 12767
rect 6837 12733 6871 12767
rect 2053 12597 2087 12631
rect 4813 12597 4847 12631
rect 8953 12597 8987 12631
rect 6745 12393 6779 12427
rect 8033 12257 8067 12291
rect 3249 12189 3283 12223
rect 3801 12189 3835 12223
rect 4445 12189 4479 12223
rect 4813 12189 4847 12223
rect 6285 12189 6319 12223
rect 8953 12189 8987 12223
rect 9137 12189 9171 12223
rect 2973 12121 3007 12155
rect 1501 12053 1535 12087
rect 3893 12053 3927 12087
rect 7481 12053 7515 12087
rect 9321 12053 9355 12087
rect 8125 11849 8159 11883
rect 9137 11849 9171 11883
rect 5825 11781 5859 11815
rect 8953 11713 8987 11747
rect 9229 11713 9263 11747
rect 3341 11645 3375 11679
rect 3617 11645 3651 11679
rect 6377 11645 6411 11679
rect 6653 11645 6687 11679
rect 1869 11509 1903 11543
rect 4353 11509 4387 11543
rect 8769 11509 8803 11543
rect 3249 11305 3283 11339
rect 8217 11237 8251 11271
rect 9137 11237 9171 11271
rect 4353 11169 4387 11203
rect 4997 11169 5031 11203
rect 1593 11101 1627 11135
rect 2605 11101 2639 11135
rect 7205 11101 7239 11135
rect 8401 11101 8435 11135
rect 8953 11101 8987 11135
rect 2145 11033 2179 11067
rect 5549 11033 5583 11067
rect 8125 11033 8159 11067
rect 8309 11033 8343 11067
rect 5825 10761 5859 10795
rect 2053 10693 2087 10727
rect 5457 10693 5491 10727
rect 1869 10625 1903 10659
rect 2881 10625 2915 10659
rect 4353 10625 4387 10659
rect 5641 10625 5675 10659
rect 6745 10625 6779 10659
rect 8217 10625 8251 10659
rect 9321 10625 9355 10659
rect 2513 10557 2547 10591
rect 6377 10557 6411 10591
rect 8677 10489 8711 10523
rect 1685 10421 1719 10455
rect 4813 10421 4847 10455
rect 9137 10421 9171 10455
rect 8953 10217 8987 10251
rect 9137 10217 9171 10251
rect 4077 10081 4111 10115
rect 6009 10081 6043 10115
rect 8309 10081 8343 10115
rect 1593 10013 1627 10047
rect 1777 10013 1811 10047
rect 2513 10013 2547 10047
rect 3801 10013 3835 10047
rect 6377 10013 6411 10047
rect 7849 10013 7883 10047
rect 9321 9945 9355 9979
rect 1961 9877 1995 9911
rect 3065 9877 3099 9911
rect 5549 9877 5583 9911
rect 8033 9877 8067 9911
rect 9121 9877 9155 9911
rect 1593 9605 1627 9639
rect 7389 9605 7423 9639
rect 9137 9605 9171 9639
rect 1777 9537 1811 9571
rect 2421 9537 2455 9571
rect 3525 9537 3559 9571
rect 5365 9537 5399 9571
rect 6469 9537 6503 9571
rect 3893 9469 3927 9503
rect 5825 9469 5859 9503
rect 1961 9333 1995 9367
rect 3065 9333 3099 9367
rect 6745 9333 6779 9367
rect 6929 9333 6963 9367
rect 1758 9129 1792 9163
rect 3249 9129 3283 9163
rect 4721 9129 4755 9163
rect 1501 8993 1535 9027
rect 4077 8993 4111 9027
rect 5273 8925 5307 8959
rect 7481 8925 7515 8959
rect 9045 8925 9079 8959
rect 7757 8857 7791 8891
rect 6561 8789 6595 8823
rect 9137 8789 9171 8823
rect 6377 8585 6411 8619
rect 9137 8517 9171 8551
rect 1961 8449 1995 8483
rect 2789 8449 2823 8483
rect 4629 8449 4663 8483
rect 5549 8449 5583 8483
rect 6929 8449 6963 8483
rect 3157 8381 3191 8415
rect 5089 8381 5123 8415
rect 8217 8381 8251 8415
rect 9321 8381 9355 8415
rect 1777 8313 1811 8347
rect 5733 8313 5767 8347
rect 1961 8041 1995 8075
rect 3801 8041 3835 8075
rect 3249 7837 3283 7871
rect 4353 7837 4387 7871
rect 7021 7837 7055 7871
rect 8033 7837 8067 7871
rect 8953 7837 8987 7871
rect 9137 7769 9171 7803
rect 5733 7701 5767 7735
rect 7481 7701 7515 7735
rect 9321 7701 9355 7735
rect 5825 7497 5859 7531
rect 9137 7497 9171 7531
rect 3617 7429 3651 7463
rect 2053 7361 2087 7395
rect 8217 7361 8251 7395
rect 9321 7361 9355 7395
rect 4077 7293 4111 7327
rect 4353 7293 4387 7327
rect 6377 7293 6411 7327
rect 6745 7293 6779 7327
rect 8677 7225 8711 7259
rect 1764 6953 1798 6987
rect 1501 6817 1535 6851
rect 3249 6817 3283 6851
rect 3893 6817 3927 6851
rect 5641 6749 5675 6783
rect 6101 6749 6135 6783
rect 6469 6749 6503 6783
rect 7941 6749 7975 6783
rect 9321 6749 9355 6783
rect 5365 6681 5399 6715
rect 8953 6681 8987 6715
rect 9137 6681 9171 6715
rect 8401 6613 8435 6647
rect 2237 6409 2271 6443
rect 3341 6409 3375 6443
rect 5733 6409 5767 6443
rect 4813 6341 4847 6375
rect 1685 6273 1719 6307
rect 2421 6273 2455 6307
rect 5549 6273 5583 6307
rect 7021 6273 7055 6307
rect 8493 6273 8527 6307
rect 5089 6205 5123 6239
rect 6653 6205 6687 6239
rect 1501 6137 1535 6171
rect 8953 6069 8987 6103
rect 2881 5865 2915 5899
rect 5549 5865 5583 5899
rect 9137 5865 9171 5899
rect 1501 5797 1535 5831
rect 2237 5729 2271 5763
rect 3801 5729 3835 5763
rect 6837 5729 6871 5763
rect 8217 5729 8251 5763
rect 1409 5661 1443 5695
rect 2145 5661 2179 5695
rect 2329 5661 2363 5695
rect 2973 5661 3007 5695
rect 8125 5661 8159 5695
rect 8953 5661 8987 5695
rect 4077 5593 4111 5627
rect 3893 5321 3927 5355
rect 4629 5321 4663 5355
rect 5733 5321 5767 5355
rect 6837 5321 6871 5355
rect 7297 5253 7331 5287
rect 9229 5253 9263 5287
rect 3801 5185 3835 5219
rect 3985 5185 4019 5219
rect 4445 5185 4479 5219
rect 4629 5185 4663 5219
rect 6193 5185 6227 5219
rect 7481 5185 7515 5219
rect 8953 5185 8987 5219
rect 9045 5185 9079 5219
rect 5089 5117 5123 5151
rect 7665 4981 7699 5015
rect 8953 4981 8987 5015
rect 6009 4777 6043 4811
rect 6745 4777 6779 4811
rect 7389 4777 7423 4811
rect 8401 4777 8435 4811
rect 4905 4641 4939 4675
rect 3525 4573 3559 4607
rect 3709 4573 3743 4607
rect 4353 4573 4387 4607
rect 6193 4573 6227 4607
rect 6837 4573 6871 4607
rect 7297 4573 7331 4607
rect 8585 4573 8619 4607
rect 9229 4573 9263 4607
rect 9321 4505 9355 4539
rect 3709 4437 3743 4471
rect 4905 4233 4939 4267
rect 3709 4097 3743 4131
rect 4997 4097 5031 4131
rect 5457 4097 5491 4131
rect 6101 4097 6135 4131
rect 6929 4097 6963 4131
rect 7849 4097 7883 4131
rect 9045 4097 9079 4131
rect 4077 4029 4111 4063
rect 6837 4029 6871 4063
rect 6285 3961 6319 3995
rect 5549 3893 5583 3927
rect 7757 3893 7791 3927
rect 9229 3893 9263 3927
rect 3709 3689 3743 3723
rect 4261 3689 4295 3723
rect 4905 3689 4939 3723
rect 6101 3689 6135 3723
rect 6837 3689 6871 3723
rect 7481 3689 7515 3723
rect 8033 3689 8067 3723
rect 3525 3485 3559 3519
rect 4169 3485 4203 3519
rect 4353 3485 4387 3519
rect 4813 3485 4847 3519
rect 4997 3485 5031 3519
rect 5917 3485 5951 3519
rect 6745 3485 6779 3519
rect 6929 3485 6963 3519
rect 7389 3485 7423 3519
rect 7573 3485 7607 3519
rect 8217 3485 8251 3519
rect 9045 3485 9079 3519
rect 9229 3349 9263 3383
rect 3709 3145 3743 3179
rect 4997 3145 5031 3179
rect 5733 3145 5767 3179
rect 6193 3145 6227 3179
rect 6929 3145 6963 3179
rect 7941 3145 7975 3179
rect 9229 3145 9263 3179
rect 3525 3009 3559 3043
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 4905 3009 4939 3043
rect 5549 3009 5583 3043
rect 5733 3009 5767 3043
rect 6377 3009 6411 3043
rect 6837 3009 6871 3043
rect 7757 3009 7791 3043
rect 9045 3009 9079 3043
rect 4169 2805 4203 2839
rect 4261 2601 4295 2635
rect 6561 2601 6595 2635
rect 8493 2601 8527 2635
rect 3709 2397 3743 2431
rect 4169 2397 4203 2431
rect 4813 2397 4847 2431
rect 4997 2397 5031 2431
rect 5917 2397 5951 2431
rect 6745 2397 6779 2431
rect 8401 2397 8435 2431
rect 8585 2397 8619 2431
rect 9229 2397 9263 2431
rect 3617 2261 3651 2295
rect 4905 2261 4939 2295
rect 6009 2261 6043 2295
rect 9045 2261 9079 2295
rect 3617 2057 3651 2091
rect 5641 2057 5675 2091
rect 8585 2057 8619 2091
rect 9229 2057 9263 2091
rect 4905 1989 4939 2023
rect 3525 1921 3559 1955
rect 3709 1921 3743 1955
rect 4169 1921 4203 1955
rect 4813 1921 4847 1955
rect 4997 1921 5031 1955
rect 5457 1921 5491 1955
rect 5641 1921 5675 1955
rect 6101 1921 6135 1955
rect 6745 1921 6779 1955
rect 6929 1921 6963 1955
rect 8677 1921 8711 1955
rect 9321 1921 9355 1955
rect 4261 1785 4295 1819
rect 6285 1717 6319 1751
rect 6837 1717 6871 1751
rect 8953 1445 8987 1479
rect 3525 1309 3559 1343
rect 4353 1309 4387 1343
rect 4813 1309 4847 1343
rect 4997 1309 5031 1343
rect 5917 1309 5951 1343
rect 6101 1309 6135 1343
rect 6745 1309 6779 1343
rect 7205 1309 7239 1343
rect 7389 1309 7423 1343
rect 4261 1241 4295 1275
rect 3709 1173 3743 1207
rect 4997 1173 5031 1207
rect 6101 1173 6135 1207
rect 6561 1173 6595 1207
rect 7389 1173 7423 1207
rect 9137 1173 9171 1207
<< metal1 >>
rect 3234 15852 3240 15904
rect 3292 15892 3298 15904
rect 8478 15892 8484 15904
rect 3292 15864 8484 15892
rect 3292 15852 3298 15864
rect 8478 15852 8484 15864
rect 8536 15852 8542 15904
rect 920 15802 9844 15824
rect 920 15750 2566 15802
rect 2618 15750 2630 15802
rect 2682 15750 2694 15802
rect 2746 15750 2758 15802
rect 2810 15750 2822 15802
rect 2874 15750 7566 15802
rect 7618 15750 7630 15802
rect 7682 15750 7694 15802
rect 7746 15750 7758 15802
rect 7810 15750 7822 15802
rect 7874 15750 9844 15802
rect 920 15728 9844 15750
rect 3237 15691 3295 15697
rect 3237 15657 3249 15691
rect 3283 15688 3295 15691
rect 4062 15688 4068 15700
rect 3283 15660 4068 15688
rect 3283 15657 3295 15660
rect 3237 15651 3295 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 9122 15688 9128 15700
rect 9083 15660 9128 15688
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 5442 15552 5448 15564
rect 5403 15524 5448 15552
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 8110 15552 8116 15564
rect 8071 15524 8116 15552
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 2682 15484 2688 15496
rect 1811 15456 2688 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 4062 15484 4068 15496
rect 4023 15456 4068 15484
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 5718 15484 5724 15496
rect 5679 15456 5724 15484
rect 5718 15444 5724 15456
rect 5776 15444 5782 15496
rect 8386 15444 8392 15496
rect 8444 15484 8450 15496
rect 8941 15487 8999 15493
rect 8444 15456 8489 15484
rect 8444 15444 8450 15456
rect 8941 15453 8953 15487
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 1394 15376 1400 15428
rect 1452 15416 1458 15428
rect 2130 15416 2136 15428
rect 1452 15388 2136 15416
rect 1452 15376 1458 15388
rect 2130 15376 2136 15388
rect 2188 15416 2194 15428
rect 2869 15419 2927 15425
rect 2869 15416 2881 15419
rect 2188 15388 2881 15416
rect 2188 15376 2194 15388
rect 2869 15385 2881 15388
rect 2915 15385 2927 15419
rect 2869 15379 2927 15385
rect 3053 15419 3111 15425
rect 3053 15385 3065 15419
rect 3099 15416 3111 15419
rect 3142 15416 3148 15428
rect 3099 15388 3148 15416
rect 3099 15385 3111 15388
rect 3053 15379 3111 15385
rect 3142 15376 3148 15388
rect 3200 15376 3206 15428
rect 4614 15416 4620 15428
rect 4575 15388 4620 15416
rect 4614 15376 4620 15388
rect 4672 15376 4678 15428
rect 7374 15376 7380 15428
rect 7432 15376 7438 15428
rect 8018 15376 8024 15428
rect 8076 15416 8082 15428
rect 8956 15416 8984 15447
rect 8076 15388 8984 15416
rect 8076 15376 8082 15388
rect 16666 15376 16672 15428
rect 16724 15376 16730 15428
rect 1210 15308 1216 15360
rect 1268 15348 1274 15360
rect 1581 15351 1639 15357
rect 1581 15348 1593 15351
rect 1268 15320 1593 15348
rect 1268 15308 1274 15320
rect 1581 15317 1593 15320
rect 1627 15317 1639 15351
rect 1581 15311 1639 15317
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 6641 15351 6699 15357
rect 6641 15348 6653 15351
rect 5592 15320 6653 15348
rect 5592 15308 5598 15320
rect 6641 15317 6653 15320
rect 6687 15317 6699 15351
rect 6641 15311 6699 15317
rect 920 15258 9844 15280
rect 920 15206 3566 15258
rect 3618 15206 3630 15258
rect 3682 15206 3694 15258
rect 3746 15206 3758 15258
rect 3810 15206 3822 15258
rect 3874 15206 8566 15258
rect 8618 15206 8630 15258
rect 8682 15206 8694 15258
rect 8746 15206 8758 15258
rect 8810 15206 8822 15258
rect 8874 15206 9844 15258
rect 920 15184 9844 15206
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 6641 15147 6699 15153
rect 6641 15144 6653 15147
rect 5776 15116 6653 15144
rect 5776 15104 5782 15116
rect 6641 15113 6653 15116
rect 6687 15113 6699 15147
rect 6641 15107 6699 15113
rect 15378 15104 15384 15156
rect 15436 15144 15442 15156
rect 16574 15144 16580 15156
rect 15436 15116 16580 15144
rect 15436 15104 15442 15116
rect 16574 15104 16580 15116
rect 16632 15104 16638 15156
rect 474 15036 480 15088
rect 532 15076 538 15088
rect 2041 15079 2099 15085
rect 2041 15076 2053 15079
rect 532 15048 2053 15076
rect 532 15036 538 15048
rect 2041 15045 2053 15048
rect 2087 15045 2099 15079
rect 2041 15039 2099 15045
rect 3237 15079 3295 15085
rect 3237 15045 3249 15079
rect 3283 15076 3295 15079
rect 4062 15076 4068 15088
rect 3283 15048 4068 15076
rect 3283 15045 3295 15048
rect 3237 15039 3295 15045
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 7374 15036 7380 15088
rect 7432 15036 7438 15088
rect 8113 15079 8171 15085
rect 8113 15045 8125 15079
rect 8159 15076 8171 15079
rect 8202 15076 8208 15088
rect 8159 15048 8208 15076
rect 8159 15045 8171 15048
rect 8113 15039 8171 15045
rect 8202 15036 8208 15048
rect 8260 15036 8266 15088
rect 1397 15011 1455 15017
rect 1397 14977 1409 15011
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 15008 2283 15011
rect 3053 15011 3111 15017
rect 3053 15008 3065 15011
rect 2271 14980 3065 15008
rect 2271 14977 2283 14980
rect 2225 14971 2283 14977
rect 3053 14977 3065 14980
rect 3099 15008 3111 15011
rect 3142 15008 3148 15020
rect 3099 14980 3148 15008
rect 3099 14977 3111 14980
rect 3053 14971 3111 14977
rect 1412 14940 1440 14971
rect 3142 14968 3148 14980
rect 3200 14968 3206 15020
rect 9033 15011 9091 15017
rect 9033 14977 9045 15011
rect 9079 15008 9091 15011
rect 9858 15008 9864 15020
rect 9079 14980 9864 15008
rect 9079 14977 9091 14980
rect 9033 14971 9091 14977
rect 9858 14968 9864 14980
rect 9916 14968 9922 15020
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 16684 15008 16712 15376
rect 16632 14980 16712 15008
rect 16632 14968 16638 14980
rect 2958 14940 2964 14952
rect 1412 14912 2964 14940
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14940 3847 14943
rect 4246 14940 4252 14952
rect 3835 14912 4252 14940
rect 3835 14909 3847 14912
rect 3789 14903 3847 14909
rect 4246 14900 4252 14912
rect 4304 14900 4310 14952
rect 4338 14900 4344 14952
rect 4396 14940 4402 14952
rect 5350 14940 5356 14952
rect 4396 14912 4441 14940
rect 5311 14912 5356 14940
rect 4396 14900 4402 14912
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 8386 14940 8392 14952
rect 8347 14912 8392 14940
rect 8386 14900 8392 14912
rect 8444 14900 8450 14952
rect 290 14832 296 14884
rect 348 14872 354 14884
rect 2409 14875 2467 14881
rect 2409 14872 2421 14875
rect 348 14844 2421 14872
rect 348 14832 354 14844
rect 2409 14841 2421 14844
rect 2455 14841 2467 14875
rect 2409 14835 2467 14841
rect 2774 14832 2780 14884
rect 2832 14872 2838 14884
rect 3234 14872 3240 14884
rect 2832 14844 3240 14872
rect 2832 14832 2838 14844
rect 3234 14832 3240 14844
rect 3292 14832 3298 14884
rect 4798 14872 4804 14884
rect 4759 14844 4804 14872
rect 4798 14832 4804 14844
rect 4856 14832 4862 14884
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 2869 14807 2927 14813
rect 2869 14773 2881 14807
rect 2915 14804 2927 14807
rect 3878 14804 3884 14816
rect 2915 14776 3884 14804
rect 2915 14773 2927 14776
rect 2869 14767 2927 14773
rect 3878 14764 3884 14776
rect 3936 14764 3942 14816
rect 9214 14804 9220 14816
rect 9175 14776 9220 14804
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 920 14714 9844 14736
rect 920 14662 2566 14714
rect 2618 14662 2630 14714
rect 2682 14662 2694 14714
rect 2746 14662 2758 14714
rect 2810 14662 2822 14714
rect 2874 14662 7566 14714
rect 7618 14662 7630 14714
rect 7682 14662 7694 14714
rect 7746 14662 7758 14714
rect 7810 14662 7822 14714
rect 7874 14662 9844 14714
rect 920 14640 9844 14662
rect 750 14560 756 14612
rect 808 14600 814 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 808 14572 4169 14600
rect 808 14560 814 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 4157 14563 4215 14569
rect 3234 14464 3240 14476
rect 3147 14436 3240 14464
rect 3234 14424 3240 14436
rect 3292 14464 3298 14476
rect 4062 14464 4068 14476
rect 3292 14436 4068 14464
rect 3292 14424 3298 14436
rect 4062 14424 4068 14436
rect 4120 14424 4126 14476
rect 4801 14467 4859 14473
rect 4801 14433 4813 14467
rect 4847 14464 4859 14467
rect 5442 14464 5448 14476
rect 4847 14436 5448 14464
rect 4847 14433 4859 14436
rect 4801 14427 4859 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 8202 14396 8208 14408
rect 8159 14368 8208 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 2498 14288 2504 14340
rect 2556 14288 2562 14340
rect 2961 14331 3019 14337
rect 2961 14297 2973 14331
rect 3007 14328 3019 14331
rect 5350 14328 5356 14340
rect 3007 14300 5356 14328
rect 3007 14297 3019 14300
rect 2961 14291 3019 14297
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 7006 14328 7012 14340
rect 6967 14300 7012 14328
rect 7006 14288 7012 14300
rect 7064 14288 7070 14340
rect 8386 14288 8392 14340
rect 8444 14328 8450 14340
rect 8941 14331 8999 14337
rect 8941 14328 8953 14331
rect 8444 14300 8953 14328
rect 8444 14288 8450 14300
rect 8941 14297 8953 14300
rect 8987 14297 8999 14331
rect 8941 14291 8999 14297
rect 9125 14331 9183 14337
rect 9125 14297 9137 14331
rect 9171 14328 9183 14331
rect 9214 14328 9220 14340
rect 9171 14300 9220 14328
rect 9171 14297 9183 14300
rect 9125 14291 9183 14297
rect 9214 14288 9220 14300
rect 9272 14288 9278 14340
rect 1489 14263 1547 14269
rect 1489 14229 1501 14263
rect 1535 14260 1547 14263
rect 1578 14260 1584 14272
rect 1535 14232 1584 14260
rect 1535 14229 1547 14232
rect 1489 14223 1547 14229
rect 1578 14220 1584 14232
rect 1636 14220 1642 14272
rect 3142 14220 3148 14272
rect 3200 14260 3206 14272
rect 4062 14260 4068 14272
rect 3200 14232 4068 14260
rect 3200 14220 3206 14232
rect 4062 14220 4068 14232
rect 4120 14220 4126 14272
rect 5534 14260 5540 14272
rect 5495 14232 5540 14260
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 7098 14220 7104 14272
rect 7156 14260 7162 14272
rect 7469 14263 7527 14269
rect 7469 14260 7481 14263
rect 7156 14232 7481 14260
rect 7156 14220 7162 14232
rect 7469 14229 7481 14232
rect 7515 14229 7527 14263
rect 9306 14260 9312 14272
rect 9267 14232 9312 14260
rect 7469 14223 7527 14229
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 920 14170 9844 14192
rect 920 14118 3566 14170
rect 3618 14118 3630 14170
rect 3682 14118 3694 14170
rect 3746 14118 3758 14170
rect 3810 14118 3822 14170
rect 3874 14118 8566 14170
rect 8618 14118 8630 14170
rect 8682 14118 8694 14170
rect 8746 14118 8758 14170
rect 8810 14118 8822 14170
rect 8874 14118 9844 14170
rect 920 14096 9844 14118
rect 3602 14016 3608 14068
rect 3660 14056 3666 14068
rect 4798 14056 4804 14068
rect 3660 14028 4804 14056
rect 3660 14016 3666 14028
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5718 14056 5724 14068
rect 5679 14028 5724 14056
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 9214 14056 9220 14068
rect 5828 14028 9220 14056
rect 3326 13948 3332 14000
rect 3384 13948 3390 14000
rect 5258 13948 5264 14000
rect 5316 13988 5322 14000
rect 5537 13991 5595 13997
rect 5537 13988 5549 13991
rect 5316 13960 5549 13988
rect 5316 13948 5322 13960
rect 5537 13957 5549 13960
rect 5583 13988 5595 13991
rect 5828 13988 5856 14028
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 5583 13960 5856 13988
rect 5583 13957 5595 13960
rect 5537 13951 5595 13957
rect 8110 13948 8116 14000
rect 8168 13948 8174 14000
rect 1302 13880 1308 13932
rect 1360 13920 1366 13932
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 1360 13892 2605 13920
rect 1360 13880 1366 13892
rect 2593 13889 2605 13892
rect 2639 13889 2651 13923
rect 4430 13920 4436 13932
rect 4391 13892 4436 13920
rect 2593 13883 2651 13889
rect 4430 13880 4436 13892
rect 4488 13880 4494 13932
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13889 5411 13923
rect 6638 13920 6644 13932
rect 6599 13892 6644 13920
rect 5353 13883 5411 13889
rect 1578 13852 1584 13864
rect 1491 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13852 1642 13864
rect 2038 13852 2044 13864
rect 1636 13824 2044 13852
rect 1636 13812 1642 13824
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 2406 13852 2412 13864
rect 2179 13824 2412 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 2406 13812 2412 13824
rect 2464 13812 2470 13864
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13852 3019 13855
rect 3602 13852 3608 13864
rect 3007 13824 3608 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 4890 13852 4896 13864
rect 4851 13824 4896 13852
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 4706 13744 4712 13796
rect 4764 13784 4770 13796
rect 5368 13784 5396 13883
rect 6638 13880 6644 13892
rect 6696 13880 6702 13932
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13920 7067 13923
rect 7098 13920 7104 13932
rect 7055 13892 7104 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13920 8539 13923
rect 9582 13920 9588 13932
rect 8527 13892 9588 13920
rect 8527 13889 8539 13892
rect 8481 13883 8539 13889
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 8938 13852 8944 13864
rect 8899 13824 8944 13852
rect 8938 13812 8944 13824
rect 8996 13812 9002 13864
rect 4764 13756 5396 13784
rect 4764 13744 4770 13756
rect 920 13626 9844 13648
rect 920 13574 2566 13626
rect 2618 13574 2630 13626
rect 2682 13574 2694 13626
rect 2746 13574 2758 13626
rect 2810 13574 2822 13626
rect 2874 13574 7566 13626
rect 7618 13574 7630 13626
rect 7682 13574 7694 13626
rect 7746 13574 7758 13626
rect 7810 13574 7822 13626
rect 7874 13574 9844 13626
rect 920 13552 9844 13574
rect 7469 13515 7527 13521
rect 7469 13481 7481 13515
rect 7515 13512 7527 13515
rect 8018 13512 8024 13524
rect 7515 13484 8024 13512
rect 7515 13481 7527 13484
rect 7469 13475 7527 13481
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 4433 13379 4491 13385
rect 4433 13376 4445 13379
rect 4212 13348 4445 13376
rect 4212 13336 4218 13348
rect 4433 13345 4445 13348
rect 4479 13376 4491 13379
rect 5258 13376 5264 13388
rect 4479 13348 5264 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 5537 13379 5595 13385
rect 5537 13345 5549 13379
rect 5583 13376 5595 13379
rect 5718 13376 5724 13388
rect 5583 13348 5724 13376
rect 5583 13345 5595 13348
rect 5537 13339 5595 13345
rect 5718 13336 5724 13348
rect 5776 13336 5782 13388
rect 16114 13336 16120 13388
rect 16172 13376 16178 13388
rect 16666 13376 16672 13388
rect 16172 13348 16672 13376
rect 16172 13336 16178 13348
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 3234 13268 3240 13320
rect 3292 13308 3298 13320
rect 3881 13311 3939 13317
rect 3881 13308 3893 13311
rect 3292 13280 3893 13308
rect 3292 13268 3298 13280
rect 3881 13277 3893 13280
rect 3927 13277 3939 13311
rect 5166 13308 5172 13320
rect 5127 13280 5172 13308
rect 3881 13271 3939 13277
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 7926 13308 7932 13320
rect 7055 13280 7932 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13277 8079 13311
rect 8938 13308 8944 13320
rect 8899 13280 8944 13308
rect 8021 13271 8079 13277
rect 1489 13243 1547 13249
rect 1489 13209 1501 13243
rect 1535 13240 1547 13243
rect 2314 13240 2320 13252
rect 1535 13212 2320 13240
rect 1535 13209 1547 13212
rect 1489 13203 1547 13209
rect 2314 13200 2320 13212
rect 2372 13200 2378 13252
rect 6638 13200 6644 13252
rect 6696 13200 6702 13252
rect 6914 13200 6920 13252
rect 6972 13240 6978 13252
rect 8036 13240 8064 13271
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 10134 13268 10140 13320
rect 10192 13308 10198 13320
rect 14274 13308 14280 13320
rect 10192 13280 14280 13308
rect 10192 13268 10198 13280
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 6972 13212 8064 13240
rect 6972 13200 6978 13212
rect 934 13132 940 13184
rect 992 13172 998 13184
rect 2777 13175 2835 13181
rect 2777 13172 2789 13175
rect 992 13144 2789 13172
rect 992 13132 998 13144
rect 2777 13141 2789 13144
rect 2823 13141 2835 13175
rect 8202 13172 8208 13184
rect 8163 13144 8208 13172
rect 2777 13135 2835 13141
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 9122 13172 9128 13184
rect 9083 13144 9128 13172
rect 9122 13132 9128 13144
rect 9180 13132 9186 13184
rect 920 13082 9844 13104
rect 920 13030 3566 13082
rect 3618 13030 3630 13082
rect 3682 13030 3694 13082
rect 3746 13030 3758 13082
rect 3810 13030 3822 13082
rect 3874 13030 8566 13082
rect 8618 13030 8630 13082
rect 8682 13030 8694 13082
rect 8746 13030 8758 13082
rect 8810 13030 8822 13082
rect 8874 13030 9844 13082
rect 920 13008 9844 13030
rect 8294 12968 8300 12980
rect 8255 12940 8300 12968
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 10318 12928 10324 12980
rect 10376 12968 10382 12980
rect 15746 12968 15752 12980
rect 10376 12940 15752 12968
rect 10376 12928 10382 12940
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 3878 12860 3884 12912
rect 3936 12860 3942 12912
rect 7282 12860 7288 12912
rect 7340 12860 7346 12912
rect 1489 12835 1547 12841
rect 1489 12801 1501 12835
rect 1535 12832 1547 12835
rect 1578 12832 1584 12844
rect 1535 12804 1584 12832
rect 1535 12801 1547 12804
rect 1489 12795 1547 12801
rect 1578 12792 1584 12804
rect 1636 12792 1642 12844
rect 2406 12792 2412 12844
rect 2464 12832 2470 12844
rect 2869 12835 2927 12841
rect 2869 12832 2881 12835
rect 2464 12804 2881 12832
rect 2464 12792 2470 12804
rect 2869 12801 2881 12804
rect 2915 12801 2927 12835
rect 4338 12832 4344 12844
rect 4299 12804 4344 12832
rect 2869 12795 2927 12801
rect 4338 12792 4344 12804
rect 4396 12792 4402 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5442 12832 5448 12844
rect 5399 12804 5448 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 9214 12832 9220 12844
rect 9175 12804 9220 12832
rect 9214 12792 9220 12804
rect 9272 12792 9278 12844
rect 2498 12764 2504 12776
rect 2459 12736 2504 12764
rect 2498 12724 2504 12736
rect 2556 12724 2562 12776
rect 5629 12767 5687 12773
rect 5629 12733 5641 12767
rect 5675 12764 5687 12767
rect 5810 12764 5816 12776
rect 5675 12736 5816 12764
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 5810 12724 5816 12736
rect 5868 12724 5874 12776
rect 6362 12724 6368 12776
rect 6420 12764 6426 12776
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 6420 12736 6561 12764
rect 6420 12724 6426 12736
rect 6549 12733 6561 12736
rect 6595 12733 6607 12767
rect 6549 12727 6607 12733
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 7190 12764 7196 12776
rect 6871 12736 7196 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 16022 12764 16028 12776
rect 10008 12736 16028 12764
rect 10008 12724 10014 12736
rect 16022 12724 16028 12736
rect 16080 12724 16086 12776
rect 106 12588 112 12640
rect 164 12628 170 12640
rect 2041 12631 2099 12637
rect 2041 12628 2053 12631
rect 164 12600 2053 12628
rect 164 12588 170 12600
rect 2041 12597 2053 12600
rect 2087 12597 2099 12631
rect 4798 12628 4804 12640
rect 4759 12600 4804 12628
rect 2041 12591 2099 12597
rect 4798 12588 4804 12600
rect 4856 12588 4862 12640
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 7926 12628 7932 12640
rect 7340 12600 7932 12628
rect 7340 12588 7346 12600
rect 7926 12588 7932 12600
rect 7984 12628 7990 12640
rect 8941 12631 8999 12637
rect 8941 12628 8953 12631
rect 7984 12600 8953 12628
rect 7984 12588 7990 12600
rect 8941 12597 8953 12600
rect 8987 12628 8999 12631
rect 9582 12628 9588 12640
rect 8987 12600 9588 12628
rect 8987 12597 8999 12600
rect 8941 12591 8999 12597
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 920 12538 9844 12560
rect 920 12486 2566 12538
rect 2618 12486 2630 12538
rect 2682 12486 2694 12538
rect 2746 12486 2758 12538
rect 2810 12486 2822 12538
rect 2874 12486 7566 12538
rect 7618 12486 7630 12538
rect 7682 12486 7694 12538
rect 7746 12486 7758 12538
rect 7810 12486 7822 12538
rect 7874 12486 9844 12538
rect 920 12464 9844 12486
rect 6733 12427 6791 12433
rect 6733 12393 6745 12427
rect 6779 12424 6791 12427
rect 6822 12424 6828 12436
rect 6779 12396 6828 12424
rect 6779 12393 6791 12396
rect 6733 12387 6791 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 9122 12384 9128 12436
rect 9180 12424 9186 12436
rect 16390 12424 16396 12436
rect 9180 12396 16396 12424
rect 9180 12384 9186 12396
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 13814 12316 13820 12368
rect 13872 12356 13878 12368
rect 14274 12356 14280 12368
rect 13872 12328 14280 12356
rect 13872 12316 13878 12328
rect 14274 12316 14280 12328
rect 14332 12316 14338 12368
rect 2958 12248 2964 12300
rect 3016 12288 3022 12300
rect 3016 12260 3832 12288
rect 3016 12248 3022 12260
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12220 3295 12223
rect 3326 12220 3332 12232
rect 3283 12192 3332 12220
rect 3283 12189 3295 12192
rect 3237 12183 3295 12189
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 3804 12229 3832 12260
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 8021 12291 8079 12297
rect 8021 12288 8033 12291
rect 7248 12260 8033 12288
rect 7248 12248 7254 12260
rect 8021 12257 8033 12260
rect 8067 12288 8079 12291
rect 8110 12288 8116 12300
rect 8067 12260 8116 12288
rect 8067 12257 8079 12260
rect 8021 12251 8079 12257
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12189 3847 12223
rect 4430 12220 4436 12232
rect 4391 12192 4436 12220
rect 3789 12183 3847 12189
rect 4430 12180 4436 12192
rect 4488 12180 4494 12232
rect 4706 12180 4712 12232
rect 4764 12220 4770 12232
rect 4801 12223 4859 12229
rect 4801 12220 4813 12223
rect 4764 12192 4813 12220
rect 4764 12180 4770 12192
rect 4801 12189 4813 12192
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12220 6331 12223
rect 6822 12220 6828 12232
rect 6319 12192 6828 12220
rect 6319 12189 6331 12192
rect 6273 12183 6331 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 8938 12220 8944 12232
rect 8899 12192 8944 12220
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 9088 12192 9137 12220
rect 9088 12180 9094 12192
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 2682 12152 2688 12164
rect 2530 12124 2688 12152
rect 2682 12112 2688 12124
rect 2740 12112 2746 12164
rect 2961 12155 3019 12161
rect 2961 12121 2973 12155
rect 3007 12121 3019 12155
rect 2961 12115 3019 12121
rect 1489 12087 1547 12093
rect 1489 12053 1501 12087
rect 1535 12084 1547 12087
rect 1578 12084 1584 12096
rect 1535 12056 1584 12084
rect 1535 12053 1547 12056
rect 1489 12047 1547 12053
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 2976 12084 3004 12115
rect 5718 12112 5724 12164
rect 5776 12112 5782 12164
rect 2096 12056 3004 12084
rect 3881 12087 3939 12093
rect 2096 12044 2102 12056
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 4062 12084 4068 12096
rect 3927 12056 4068 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 7469 12087 7527 12093
rect 7469 12084 7481 12087
rect 6972 12056 7481 12084
rect 6972 12044 6978 12056
rect 7469 12053 7481 12056
rect 7515 12053 7527 12087
rect 7469 12047 7527 12053
rect 9309 12087 9367 12093
rect 9309 12053 9321 12087
rect 9355 12084 9367 12087
rect 9766 12084 9772 12096
rect 9355 12056 9772 12084
rect 9355 12053 9367 12056
rect 9309 12047 9367 12053
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 16206 12044 16212 12096
rect 16264 12084 16270 12096
rect 16390 12084 16396 12096
rect 16264 12056 16396 12084
rect 16264 12044 16270 12056
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 920 11994 9844 12016
rect 920 11942 3566 11994
rect 3618 11942 3630 11994
rect 3682 11942 3694 11994
rect 3746 11942 3758 11994
rect 3810 11942 3822 11994
rect 3874 11942 8566 11994
rect 8618 11942 8630 11994
rect 8682 11942 8694 11994
rect 8746 11942 8758 11994
rect 8810 11942 8822 11994
rect 8874 11942 9844 11994
rect 920 11920 9844 11942
rect 10502 11908 10508 11960
rect 10560 11948 10566 11960
rect 16206 11948 16212 11960
rect 10560 11920 16212 11948
rect 10560 11908 10566 11920
rect 16206 11908 16212 11920
rect 16264 11908 16270 11960
rect 7926 11880 7932 11892
rect 7024 11852 7932 11880
rect 2682 11772 2688 11824
rect 2740 11772 2746 11824
rect 3326 11772 3332 11824
rect 3384 11812 3390 11824
rect 5810 11812 5816 11824
rect 3384 11784 3648 11812
rect 5771 11784 5816 11812
rect 3384 11772 3390 11784
rect 3326 11676 3332 11688
rect 3287 11648 3332 11676
rect 3326 11636 3332 11648
rect 3384 11636 3390 11688
rect 3620 11685 3648 11784
rect 5810 11772 5816 11784
rect 5868 11772 5874 11824
rect 7024 11812 7052 11852
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 8110 11880 8116 11892
rect 8071 11852 8116 11880
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 9122 11880 9128 11892
rect 9083 11852 9128 11880
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 7098 11812 7104 11824
rect 7024 11784 7104 11812
rect 7098 11772 7104 11784
rect 7156 11772 7162 11824
rect 10686 11772 10692 11824
rect 10744 11812 10750 11824
rect 15838 11812 15844 11824
rect 10744 11784 15844 11812
rect 10744 11772 10750 11784
rect 15838 11772 15844 11784
rect 15896 11772 15902 11824
rect 8938 11744 8944 11756
rect 8899 11716 8944 11744
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 9214 11744 9220 11756
rect 9175 11716 9220 11744
rect 9214 11704 9220 11716
rect 9272 11704 9278 11756
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11676 3663 11679
rect 6270 11676 6276 11688
rect 3651 11648 6276 11676
rect 3651 11645 3663 11648
rect 3605 11639 3663 11645
rect 6270 11636 6276 11648
rect 6328 11676 6334 11688
rect 6365 11679 6423 11685
rect 6365 11676 6377 11679
rect 6328 11648 6377 11676
rect 6328 11636 6334 11648
rect 6365 11645 6377 11648
rect 6411 11645 6423 11679
rect 6638 11676 6644 11688
rect 6599 11648 6644 11676
rect 6365 11639 6423 11645
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 1854 11540 1860 11552
rect 1815 11512 1860 11540
rect 1854 11500 1860 11512
rect 1912 11500 1918 11552
rect 4338 11540 4344 11552
rect 4299 11512 4344 11540
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8757 11543 8815 11549
rect 8757 11540 8769 11543
rect 8352 11512 8769 11540
rect 8352 11500 8358 11512
rect 8757 11509 8769 11512
rect 8803 11509 8815 11543
rect 8757 11503 8815 11509
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 7566 11450
rect 7618 11398 7630 11450
rect 7682 11398 7694 11450
rect 7746 11398 7758 11450
rect 7810 11398 7822 11450
rect 7874 11398 9844 11450
rect 920 11376 9844 11398
rect 3237 11339 3295 11345
rect 3237 11305 3249 11339
rect 3283 11336 3295 11339
rect 3970 11336 3976 11348
rect 3283 11308 3976 11336
rect 3283 11305 3295 11308
rect 3237 11299 3295 11305
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 11146 11296 11152 11348
rect 11204 11336 11210 11348
rect 11422 11336 11428 11348
rect 11204 11308 11428 11336
rect 11204 11296 11210 11308
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 8202 11268 8208 11280
rect 8163 11240 8208 11268
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 9122 11268 9128 11280
rect 9083 11240 9128 11268
rect 9122 11228 9128 11240
rect 9180 11228 9186 11280
rect 566 11160 572 11212
rect 624 11200 630 11212
rect 4341 11203 4399 11209
rect 4341 11200 4353 11203
rect 624 11172 4353 11200
rect 624 11160 630 11172
rect 4341 11169 4353 11172
rect 4387 11169 4399 11203
rect 4982 11200 4988 11212
rect 4943 11172 4988 11200
rect 4341 11163 4399 11169
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 1578 11132 1584 11144
rect 1539 11104 1584 11132
rect 1578 11092 1584 11104
rect 1636 11092 1642 11144
rect 1854 11092 1860 11144
rect 1912 11132 1918 11144
rect 2593 11135 2651 11141
rect 2593 11132 2605 11135
rect 1912 11104 2605 11132
rect 1912 11092 1918 11104
rect 2593 11101 2605 11104
rect 2639 11132 2651 11135
rect 7190 11132 7196 11144
rect 2639 11104 2820 11132
rect 7151 11104 7196 11132
rect 2639 11101 2651 11104
rect 2593 11095 2651 11101
rect 2133 11067 2191 11073
rect 2133 11033 2145 11067
rect 2179 11064 2191 11067
rect 2682 11064 2688 11076
rect 2179 11036 2688 11064
rect 2179 11033 2191 11036
rect 2133 11027 2191 11033
rect 2682 11024 2688 11036
rect 2740 11024 2746 11076
rect 2792 10996 2820 11104
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 5534 11064 5540 11076
rect 5495 11036 5540 11064
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 8018 11064 8024 11076
rect 7340 11036 8024 11064
rect 7340 11024 7346 11036
rect 8018 11024 8024 11036
rect 8076 11064 8082 11076
rect 8113 11067 8171 11073
rect 8113 11064 8125 11067
rect 8076 11036 8125 11064
rect 8076 11024 8082 11036
rect 8113 11033 8125 11036
rect 8159 11033 8171 11067
rect 8113 11027 8171 11033
rect 8297 11067 8355 11073
rect 8297 11033 8309 11067
rect 8343 11033 8355 11067
rect 8404 11064 8432 11095
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8536 11104 8953 11132
rect 8536 11092 8542 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 16574 11092 16580 11144
rect 16632 11132 16638 11144
rect 16632 11104 16712 11132
rect 16632 11092 16638 11104
rect 9858 11064 9864 11076
rect 8404 11036 9864 11064
rect 8297 11027 8355 11033
rect 3142 10996 3148 11008
rect 2792 10968 3148 10996
rect 3142 10956 3148 10968
rect 3200 10956 3206 11008
rect 8312 10996 8340 11027
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 9214 10996 9220 11008
rect 8312 10968 9220 10996
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 16114 10956 16120 11008
rect 16172 10996 16178 11008
rect 16574 10996 16580 11008
rect 16172 10968 16580 10996
rect 16172 10956 16178 10968
rect 16574 10956 16580 10968
rect 16632 10956 16638 11008
rect 920 10906 9844 10928
rect 920 10854 3566 10906
rect 3618 10854 3630 10906
rect 3682 10854 3694 10906
rect 3746 10854 3758 10906
rect 3810 10854 3822 10906
rect 3874 10854 8566 10906
rect 8618 10854 8630 10906
rect 8682 10854 8694 10906
rect 8746 10854 8758 10906
rect 8810 10854 8822 10906
rect 8874 10854 9844 10906
rect 15102 10888 15108 10940
rect 15160 10928 15166 10940
rect 15470 10928 15476 10940
rect 15160 10900 15476 10928
rect 15160 10888 15166 10900
rect 15470 10888 15476 10900
rect 15528 10888 15534 10940
rect 16390 10888 16396 10940
rect 16448 10888 16454 10940
rect 920 10832 9844 10854
rect 5626 10792 5632 10804
rect 5460 10764 5632 10792
rect 2041 10727 2099 10733
rect 2041 10693 2053 10727
rect 2087 10724 2099 10727
rect 2222 10724 2228 10736
rect 2087 10696 2228 10724
rect 2087 10693 2099 10696
rect 2041 10687 2099 10693
rect 2222 10684 2228 10696
rect 2280 10684 2286 10736
rect 4154 10724 4160 10736
rect 4002 10696 4160 10724
rect 4154 10684 4160 10696
rect 4212 10684 4218 10736
rect 5460 10733 5488 10764
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 5859 10764 8340 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 5445 10727 5503 10733
rect 5445 10693 5457 10727
rect 5491 10693 5503 10727
rect 5445 10687 5503 10693
rect 7190 10684 7196 10736
rect 7248 10684 7254 10736
rect 1762 10616 1768 10668
rect 1820 10656 1826 10668
rect 1857 10659 1915 10665
rect 1857 10656 1869 10659
rect 1820 10628 1869 10656
rect 1820 10616 1826 10628
rect 1857 10625 1869 10628
rect 1903 10656 1915 10659
rect 2406 10656 2412 10668
rect 1903 10628 2412 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 2774 10616 2780 10668
rect 2832 10656 2838 10668
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2832 10628 2881 10656
rect 2832 10616 2838 10628
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 5350 10656 5356 10668
rect 4387 10628 5356 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5626 10656 5632 10668
rect 5587 10628 5632 10656
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 6822 10656 6828 10668
rect 6779 10628 6828 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 8202 10656 8208 10668
rect 8163 10628 8208 10656
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 8312 10656 8340 10764
rect 9309 10659 9367 10665
rect 9309 10656 9321 10659
rect 8312 10628 9321 10656
rect 9309 10625 9321 10628
rect 9355 10625 9367 10659
rect 16408 10656 16436 10888
rect 16408 10628 16620 10656
rect 9309 10619 9367 10625
rect 1026 10548 1032 10600
rect 1084 10588 1090 10600
rect 2501 10591 2559 10597
rect 2501 10588 2513 10591
rect 1084 10560 2513 10588
rect 1084 10548 1090 10560
rect 2501 10557 2513 10560
rect 2547 10557 2559 10591
rect 6362 10588 6368 10600
rect 6323 10560 6368 10588
rect 2501 10551 2559 10557
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 8018 10480 8024 10532
rect 8076 10520 8082 10532
rect 8665 10523 8723 10529
rect 8665 10520 8677 10523
rect 8076 10492 8677 10520
rect 8076 10480 8082 10492
rect 8665 10489 8677 10492
rect 8711 10489 8723 10523
rect 8665 10483 8723 10489
rect 13446 10480 13452 10532
rect 13504 10520 13510 10532
rect 14274 10520 14280 10532
rect 13504 10492 14280 10520
rect 13504 10480 13510 10492
rect 14274 10480 14280 10492
rect 14332 10480 14338 10532
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 15620 10492 16528 10520
rect 15620 10480 15626 10492
rect 1673 10455 1731 10461
rect 1673 10421 1685 10455
rect 1719 10452 1731 10455
rect 2222 10452 2228 10464
rect 1719 10424 2228 10452
rect 1719 10421 1731 10424
rect 1673 10415 1731 10421
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 5350 10452 5356 10464
rect 4847 10424 5356 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 9122 10452 9128 10464
rect 9083 10424 9128 10452
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 7566 10362
rect 7618 10310 7630 10362
rect 7682 10310 7694 10362
rect 7746 10310 7758 10362
rect 7810 10310 7822 10362
rect 7874 10310 9844 10362
rect 920 10288 9844 10310
rect 8938 10248 8944 10260
rect 8899 10220 8944 10248
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9125 10251 9183 10257
rect 9125 10217 9137 10251
rect 9171 10248 9183 10251
rect 9214 10248 9220 10260
rect 9171 10220 9220 10248
rect 9171 10217 9183 10220
rect 9125 10211 9183 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 15470 10208 15476 10260
rect 15528 10248 15534 10260
rect 16390 10248 16396 10260
rect 15528 10220 16396 10248
rect 15528 10208 15534 10220
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 16500 10180 16528 10492
rect 16408 10152 16528 10180
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 3200 10084 4077 10112
rect 3200 10072 3206 10084
rect 4065 10081 4077 10084
rect 4111 10081 4123 10115
rect 5994 10112 6000 10124
rect 5955 10084 6000 10112
rect 4065 10075 4123 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10112 8355 10115
rect 9214 10112 9220 10124
rect 8343 10084 9220 10112
rect 8343 10081 8355 10084
rect 8297 10075 8355 10081
rect 9214 10072 9220 10084
rect 9272 10072 9278 10124
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 14366 10112 14372 10124
rect 13964 10084 14372 10112
rect 13964 10072 13970 10084
rect 14366 10072 14372 10084
rect 14424 10072 14430 10124
rect 1486 10004 1492 10056
rect 1544 10044 1550 10056
rect 1581 10047 1639 10053
rect 1581 10044 1593 10047
rect 1544 10016 1593 10044
rect 1544 10004 1550 10016
rect 1581 10013 1593 10016
rect 1627 10013 1639 10047
rect 1762 10044 1768 10056
rect 1723 10016 1768 10044
rect 1581 10007 1639 10013
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10044 2559 10047
rect 2547 10016 2774 10044
rect 2547 10013 2559 10016
rect 2501 10007 2559 10013
rect 2746 9976 2774 10016
rect 3050 10004 3056 10056
rect 3108 10044 3114 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3108 10016 3801 10044
rect 3108 10004 3114 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 5166 10004 5172 10056
rect 5224 10004 5230 10056
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10044 6423 10047
rect 6454 10044 6460 10056
rect 6411 10016 6460 10044
rect 6411 10013 6423 10016
rect 6365 10007 6423 10013
rect 6454 10004 6460 10016
rect 6512 10004 6518 10056
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 9122 10044 9128 10056
rect 7883 10016 9128 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 16298 10044 16304 10056
rect 13780 10016 16304 10044
rect 13780 10004 13786 10016
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 3234 9976 3240 9988
rect 2746 9948 3240 9976
rect 3234 9936 3240 9948
rect 3292 9936 3298 9988
rect 7098 9936 7104 9988
rect 7156 9936 7162 9988
rect 9306 9976 9312 9988
rect 9267 9948 9312 9976
rect 9306 9936 9312 9948
rect 9364 9936 9370 9988
rect 16408 9976 16436 10152
rect 16482 10072 16488 10124
rect 16540 10072 16546 10124
rect 16132 9948 16436 9976
rect 1949 9911 2007 9917
rect 1949 9877 1961 9911
rect 1995 9908 2007 9911
rect 2314 9908 2320 9920
rect 1995 9880 2320 9908
rect 1995 9877 2007 9880
rect 1949 9871 2007 9877
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 3053 9911 3111 9917
rect 3053 9877 3065 9911
rect 3099 9908 3111 9911
rect 3142 9908 3148 9920
rect 3099 9880 3148 9908
rect 3099 9877 3111 9880
rect 3053 9871 3111 9877
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 5537 9911 5595 9917
rect 5537 9877 5549 9911
rect 5583 9908 5595 9911
rect 6638 9908 6644 9920
rect 5583 9880 6644 9908
rect 5583 9877 5595 9880
rect 5537 9871 5595 9877
rect 6638 9868 6644 9880
rect 6696 9908 6702 9920
rect 6822 9908 6828 9920
rect 6696 9880 6828 9908
rect 6696 9868 6702 9880
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 8018 9908 8024 9920
rect 7979 9880 8024 9908
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 9109 9911 9167 9917
rect 9109 9908 9121 9911
rect 8444 9880 9121 9908
rect 8444 9868 8450 9880
rect 9109 9877 9121 9880
rect 9155 9908 9167 9911
rect 9398 9908 9404 9920
rect 9155 9880 9404 9908
rect 9155 9877 9167 9880
rect 9109 9871 9167 9877
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 920 9818 9844 9840
rect 920 9766 3566 9818
rect 3618 9766 3630 9818
rect 3682 9766 3694 9818
rect 3746 9766 3758 9818
rect 3810 9766 3822 9818
rect 3874 9766 8566 9818
rect 8618 9766 8630 9818
rect 8682 9766 8694 9818
rect 8746 9766 8758 9818
rect 8810 9766 8822 9818
rect 8874 9766 9844 9818
rect 920 9744 9844 9766
rect 1762 9664 1768 9716
rect 1820 9664 1826 9716
rect 4890 9664 4896 9716
rect 4948 9704 4954 9716
rect 4948 9676 5580 9704
rect 4948 9664 4954 9676
rect 1581 9639 1639 9645
rect 1581 9605 1593 9639
rect 1627 9636 1639 9639
rect 1670 9636 1676 9648
rect 1627 9608 1676 9636
rect 1627 9605 1639 9608
rect 1581 9599 1639 9605
rect 1670 9596 1676 9608
rect 1728 9596 1734 9648
rect 1780 9577 1808 9664
rect 4614 9596 4620 9648
rect 4672 9596 4678 9648
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 2130 9528 2136 9580
rect 2188 9568 2194 9580
rect 2409 9571 2467 9577
rect 2409 9568 2421 9571
rect 2188 9540 2421 9568
rect 2188 9528 2194 9540
rect 2409 9537 2421 9540
rect 2455 9537 2467 9571
rect 2409 9531 2467 9537
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 3513 9571 3571 9577
rect 3513 9568 3525 9571
rect 3476 9540 3525 9568
rect 3476 9528 3482 9540
rect 3513 9537 3525 9540
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 5166 9528 5172 9580
rect 5224 9568 5230 9580
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 5224 9540 5365 9568
rect 5224 9528 5230 9540
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5552 9568 5580 9676
rect 7006 9596 7012 9648
rect 7064 9636 7070 9648
rect 7377 9639 7435 9645
rect 7377 9636 7389 9639
rect 7064 9608 7389 9636
rect 7064 9596 7070 9608
rect 7377 9605 7389 9608
rect 7423 9605 7435 9639
rect 9122 9636 9128 9648
rect 9083 9608 9128 9636
rect 7377 9599 7435 9605
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 6457 9571 6515 9577
rect 6457 9568 6469 9571
rect 5552 9540 6469 9568
rect 5353 9531 5411 9537
rect 6457 9537 6469 9540
rect 6503 9568 6515 9571
rect 6822 9568 6828 9580
rect 6503 9540 6828 9568
rect 6503 9537 6515 9540
rect 6457 9531 6515 9537
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9500 3939 9503
rect 4062 9500 4068 9512
rect 3927 9472 4068 9500
rect 3927 9469 3939 9472
rect 3881 9463 3939 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 5810 9500 5816 9512
rect 5771 9472 5816 9500
rect 5810 9460 5816 9472
rect 5868 9460 5874 9512
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 15378 9500 15384 9512
rect 13872 9472 15384 9500
rect 13872 9460 13878 9472
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 842 9324 848 9376
rect 900 9364 906 9376
rect 1949 9367 2007 9373
rect 1949 9364 1961 9367
rect 900 9336 1961 9364
rect 900 9324 906 9336
rect 1949 9333 1961 9336
rect 1995 9333 2007 9367
rect 1949 9327 2007 9333
rect 3053 9367 3111 9373
rect 3053 9333 3065 9367
rect 3099 9364 3111 9367
rect 3878 9364 3884 9376
rect 3099 9336 3884 9364
rect 3099 9333 3111 9336
rect 3053 9327 3111 9333
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 6730 9364 6736 9376
rect 6691 9336 6736 9364
rect 6730 9324 6736 9336
rect 6788 9324 6794 9376
rect 6917 9367 6975 9373
rect 6917 9333 6929 9367
rect 6963 9364 6975 9367
rect 9030 9364 9036 9376
rect 6963 9336 9036 9364
rect 6963 9333 6975 9336
rect 6917 9327 6975 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 15562 9364 15568 9376
rect 15344 9336 15568 9364
rect 15344 9324 15350 9336
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 7566 9274
rect 7618 9222 7630 9274
rect 7682 9222 7694 9274
rect 7746 9222 7758 9274
rect 7810 9222 7822 9274
rect 7874 9222 9844 9274
rect 920 9200 9844 9222
rect 15562 9188 15568 9240
rect 15620 9228 15626 9240
rect 15746 9228 15752 9240
rect 15620 9200 15752 9228
rect 15620 9188 15626 9200
rect 15746 9188 15752 9200
rect 15804 9188 15810 9240
rect 1578 9120 1584 9172
rect 1636 9160 1642 9172
rect 1746 9163 1804 9169
rect 1746 9160 1758 9163
rect 1636 9132 1758 9160
rect 1636 9120 1642 9132
rect 1746 9129 1758 9132
rect 1792 9129 1804 9163
rect 1746 9123 1804 9129
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 3234 9160 3240 9172
rect 2832 9132 3240 9160
rect 2832 9120 2838 9132
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 4706 9160 4712 9172
rect 4667 9132 4712 9160
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 2866 9052 2872 9104
rect 2924 9092 2930 9104
rect 3142 9092 3148 9104
rect 2924 9064 3148 9092
rect 2924 9052 2930 9064
rect 3142 9052 3148 9064
rect 3200 9052 3206 9104
rect 15746 9052 15752 9104
rect 15804 9092 15810 9104
rect 16132 9092 16160 9948
rect 16500 9852 16528 10072
rect 16482 9800 16488 9852
rect 16540 9800 16546 9852
rect 15804 9064 16160 9092
rect 15804 9052 15810 9064
rect 1489 9027 1547 9033
rect 1489 8993 1501 9027
rect 1535 9024 1547 9027
rect 3050 9024 3056 9036
rect 1535 8996 3056 9024
rect 1535 8993 1547 8996
rect 1489 8987 1547 8993
rect 3050 8984 3056 8996
rect 3108 8984 3114 9036
rect 3326 8984 3332 9036
rect 3384 9024 3390 9036
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 3384 8996 4077 9024
rect 3384 8984 3390 8996
rect 4065 8993 4077 8996
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 5261 8959 5319 8965
rect 5261 8956 5273 8959
rect 4212 8928 5273 8956
rect 4212 8916 4218 8928
rect 5261 8925 5273 8928
rect 5307 8956 5319 8959
rect 5442 8956 5448 8968
rect 5307 8928 5448 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 6546 8916 6552 8968
rect 6604 8956 6610 8968
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 6604 8928 7481 8956
rect 6604 8916 6610 8928
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 9030 8956 9036 8968
rect 8991 8928 9036 8956
rect 7469 8919 7527 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 15654 8956 15660 8968
rect 15436 8928 15660 8956
rect 15436 8916 15442 8928
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 3418 8888 3424 8900
rect 2990 8860 3424 8888
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 7374 8848 7380 8900
rect 7432 8888 7438 8900
rect 7745 8891 7803 8897
rect 7745 8888 7757 8891
rect 7432 8860 7757 8888
rect 7432 8848 7438 8860
rect 7745 8857 7757 8860
rect 7791 8857 7803 8891
rect 7745 8851 7803 8857
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 6270 8820 6276 8832
rect 5592 8792 6276 8820
rect 5592 8780 5598 8792
rect 6270 8780 6276 8792
rect 6328 8820 6334 8832
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 6328 8792 6561 8820
rect 6328 8780 6334 8792
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 9122 8820 9128 8832
rect 9083 8792 9128 8820
rect 6549 8783 6607 8789
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 15654 8780 15660 8832
rect 15712 8820 15718 8832
rect 16482 8820 16488 8832
rect 15712 8792 16488 8820
rect 15712 8780 15718 8792
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 920 8730 9844 8752
rect 920 8678 3566 8730
rect 3618 8678 3630 8730
rect 3682 8678 3694 8730
rect 3746 8678 3758 8730
rect 3810 8678 3822 8730
rect 3874 8678 8566 8730
rect 8618 8678 8630 8730
rect 8682 8678 8694 8730
rect 8746 8678 8758 8730
rect 8810 8678 8822 8730
rect 8874 8678 9844 8730
rect 920 8656 9844 8678
rect 16482 8644 16488 8696
rect 16540 8684 16546 8696
rect 16592 8684 16620 10628
rect 16540 8656 16620 8684
rect 16540 8644 16546 8656
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 6365 8619 6423 8625
rect 3292 8588 3464 8616
rect 3292 8576 3298 8588
rect 3436 8548 3464 8588
rect 6365 8585 6377 8619
rect 6411 8616 6423 8619
rect 6454 8616 6460 8628
rect 6411 8588 6460 8616
rect 6411 8585 6423 8588
rect 6365 8579 6423 8585
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 16574 8576 16580 8628
rect 16632 8576 16638 8628
rect 3436 8520 3542 8548
rect 4522 8508 4528 8560
rect 4580 8548 4586 8560
rect 9122 8548 9128 8560
rect 4580 8520 4660 8548
rect 9083 8520 9128 8548
rect 4580 8508 4586 8520
rect 1946 8480 1952 8492
rect 1907 8452 1952 8480
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 4632 8489 4660 8520
rect 9122 8508 9128 8520
rect 9180 8508 9186 8560
rect 16592 8548 16620 8576
rect 16408 8520 16620 8548
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8480 2835 8483
rect 4617 8483 4675 8489
rect 2823 8452 3280 8480
rect 2823 8449 2835 8452
rect 2777 8443 2835 8449
rect 2866 8372 2872 8424
rect 2924 8412 2930 8424
rect 3145 8415 3203 8421
rect 3145 8412 3157 8415
rect 2924 8384 3157 8412
rect 2924 8372 2930 8384
rect 3145 8381 3157 8384
rect 3191 8381 3203 8415
rect 3252 8412 3280 8452
rect 4617 8449 4629 8483
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 5626 8480 5632 8492
rect 5583 8452 5632 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 6914 8480 6920 8492
rect 6875 8452 6920 8480
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 15562 8440 15568 8492
rect 15620 8440 15626 8492
rect 3786 8412 3792 8424
rect 3252 8384 3792 8412
rect 3145 8375 3203 8381
rect 3786 8372 3792 8384
rect 3844 8372 3850 8424
rect 5077 8415 5135 8421
rect 5077 8381 5089 8415
rect 5123 8412 5135 8415
rect 6730 8412 6736 8424
rect 5123 8384 6736 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 6730 8372 6736 8384
rect 6788 8372 6794 8424
rect 8202 8412 8208 8424
rect 8163 8384 8208 8412
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8412 9367 8415
rect 9582 8412 9588 8424
rect 9355 8384 9588 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 1762 8344 1768 8356
rect 1723 8316 1768 8344
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 2774 8344 2780 8356
rect 2746 8304 2780 8344
rect 2832 8304 2838 8356
rect 5721 8347 5779 8353
rect 5721 8313 5733 8347
rect 5767 8344 5779 8347
rect 6822 8344 6828 8356
rect 5767 8316 6828 8344
rect 5767 8313 5779 8316
rect 5721 8307 5779 8313
rect 6822 8304 6828 8316
rect 6880 8304 6886 8356
rect 1946 8236 1952 8288
rect 2004 8276 2010 8288
rect 2746 8276 2774 8304
rect 2004 8248 2774 8276
rect 2004 8236 2010 8248
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 7566 8186
rect 7618 8134 7630 8186
rect 7682 8134 7694 8186
rect 7746 8134 7758 8186
rect 7810 8134 7822 8186
rect 7874 8134 9844 8186
rect 920 8112 9844 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2038 8072 2044 8084
rect 1995 8044 2044 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2038 8032 2044 8044
rect 2096 8072 2102 8084
rect 2958 8072 2964 8084
rect 2096 8044 2964 8072
rect 2096 8032 2102 8044
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3789 8075 3847 8081
rect 3789 8041 3801 8075
rect 3835 8072 3847 8075
rect 4062 8072 4068 8084
rect 3835 8044 4068 8072
rect 3835 8041 3847 8044
rect 3789 8035 3847 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 4246 7868 4252 7880
rect 3283 7840 4252 7868
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 4246 7828 4252 7840
rect 4304 7828 4310 7880
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 7006 7868 7012 7880
rect 4396 7840 4441 7868
rect 6967 7840 7012 7868
rect 4396 7828 4402 7840
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 8018 7868 8024 7880
rect 7979 7840 8024 7868
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8938 7868 8944 7880
rect 8899 7840 8944 7868
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 15580 7868 15608 8440
rect 16408 8208 16436 8520
rect 16574 8440 16580 8492
rect 16632 8440 16638 8492
rect 16592 8412 16620 8440
rect 16684 8424 16712 11104
rect 16546 8384 16620 8412
rect 16546 8288 16574 8384
rect 16666 8372 16672 8424
rect 16724 8372 16730 8424
rect 16482 8236 16488 8288
rect 16540 8248 16574 8288
rect 16540 8236 16546 8248
rect 16574 8208 16580 8220
rect 16408 8180 16580 8208
rect 16574 8168 16580 8180
rect 16632 8168 16638 8220
rect 15528 7840 15608 7868
rect 15528 7828 15534 7840
rect 9122 7800 9128 7812
rect 9083 7772 9128 7800
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 3694 7692 3700 7744
rect 3752 7732 3758 7744
rect 4246 7732 4252 7744
rect 3752 7704 4252 7732
rect 3752 7692 3758 7704
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 5721 7735 5779 7741
rect 5721 7701 5733 7735
rect 5767 7732 5779 7735
rect 6270 7732 6276 7744
rect 5767 7704 6276 7732
rect 5767 7701 5779 7704
rect 5721 7695 5779 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7469 7735 7527 7741
rect 7469 7732 7481 7735
rect 7064 7704 7481 7732
rect 7064 7692 7070 7704
rect 7469 7701 7481 7704
rect 7515 7701 7527 7735
rect 7469 7695 7527 7701
rect 9309 7735 9367 7741
rect 9309 7701 9321 7735
rect 9355 7732 9367 7735
rect 9398 7732 9404 7744
rect 9355 7704 9404 7732
rect 9355 7701 9367 7704
rect 9309 7695 9367 7701
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 920 7642 9844 7664
rect 920 7590 3566 7642
rect 3618 7590 3630 7642
rect 3682 7590 3694 7642
rect 3746 7590 3758 7642
rect 3810 7590 3822 7642
rect 3874 7590 8566 7642
rect 8618 7590 8630 7642
rect 8682 7590 8694 7642
rect 8746 7590 8758 7642
rect 8810 7590 8822 7642
rect 8874 7590 9844 7642
rect 920 7568 9844 7590
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 5408 7500 5825 7528
rect 5408 7488 5414 7500
rect 5813 7497 5825 7500
rect 5859 7528 5871 7531
rect 8018 7528 8024 7540
rect 5859 7500 8024 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8352 7500 9137 7528
rect 8352 7488 8358 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9125 7491 9183 7497
rect 3605 7463 3663 7469
rect 3605 7429 3617 7463
rect 3651 7460 3663 7463
rect 4062 7460 4068 7472
rect 3651 7432 4068 7460
rect 3651 7429 3663 7432
rect 3605 7423 3663 7429
rect 4062 7420 4068 7432
rect 4120 7420 4126 7472
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 4304 7432 4830 7460
rect 4304 7420 4310 7432
rect 7098 7420 7104 7472
rect 7156 7420 7162 7472
rect 1486 7352 1492 7404
rect 1544 7392 1550 7404
rect 2041 7395 2099 7401
rect 2041 7392 2053 7395
rect 1544 7364 2053 7392
rect 1544 7352 1550 7364
rect 2041 7361 2053 7364
rect 2087 7392 2099 7395
rect 3050 7392 3056 7404
rect 2087 7364 3056 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 8076 7364 8217 7392
rect 8076 7352 8082 7364
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 9766 7392 9772 7404
rect 9355 7364 9772 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 3068 7324 3096 7352
rect 4062 7324 4068 7336
rect 3068 7296 4068 7324
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 4341 7327 4399 7333
rect 4341 7324 4353 7327
rect 4172 7296 4353 7324
rect 3050 7216 3056 7268
rect 3108 7256 3114 7268
rect 3234 7256 3240 7268
rect 3108 7228 3240 7256
rect 3108 7216 3114 7228
rect 3234 7216 3240 7228
rect 3292 7216 3298 7268
rect 4172 7200 4200 7296
rect 4341 7293 4353 7296
rect 4387 7293 4399 7327
rect 6362 7324 6368 7336
rect 6323 7296 6368 7324
rect 4341 7287 4399 7293
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 6730 7324 6736 7336
rect 6691 7296 6736 7324
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 8665 7259 8723 7265
rect 8665 7225 8677 7259
rect 8711 7256 8723 7259
rect 9766 7256 9772 7268
rect 8711 7228 9772 7256
rect 8711 7225 8723 7228
rect 8665 7219 8723 7225
rect 9766 7216 9772 7228
rect 9824 7216 9830 7268
rect 16482 7216 16488 7268
rect 16540 7216 16546 7268
rect 4154 7148 4160 7200
rect 4212 7148 4218 7200
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 7566 7098
rect 7618 7046 7630 7098
rect 7682 7046 7694 7098
rect 7746 7046 7758 7098
rect 7810 7046 7822 7098
rect 7874 7046 9844 7098
rect 920 7024 9844 7046
rect 11330 7012 11336 7064
rect 11388 7052 11394 7064
rect 16022 7052 16028 7064
rect 11388 7024 16028 7052
rect 11388 7012 11394 7024
rect 16022 7012 16028 7024
rect 16080 7012 16086 7064
rect 16500 7052 16528 7216
rect 16574 7052 16580 7064
rect 16500 7024 16580 7052
rect 16574 7012 16580 7024
rect 16632 7012 16638 7064
rect 1752 6987 1810 6993
rect 1752 6953 1764 6987
rect 1798 6984 1810 6987
rect 1946 6984 1952 6996
rect 1798 6956 1952 6984
rect 1798 6953 1810 6956
rect 1752 6947 1810 6953
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 4338 6984 4344 6996
rect 3804 6956 4344 6984
rect 1486 6848 1492 6860
rect 1447 6820 1492 6848
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 3326 6848 3332 6860
rect 3283 6820 3332 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 3326 6808 3332 6820
rect 3384 6848 3390 6860
rect 3804 6848 3832 6956
rect 4338 6944 4344 6956
rect 4396 6944 4402 6996
rect 4154 6916 4160 6928
rect 4080 6888 4160 6916
rect 3384 6820 3832 6848
rect 3881 6851 3939 6857
rect 3384 6808 3390 6820
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 4080 6848 4108 6888
rect 4154 6876 4160 6888
rect 4212 6876 4218 6928
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 8938 6916 8944 6928
rect 8352 6888 8944 6916
rect 8352 6876 8358 6888
rect 8938 6876 8944 6888
rect 8996 6876 9002 6928
rect 3927 6820 4108 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 10594 6808 10600 6860
rect 10652 6848 10658 6860
rect 15838 6848 15844 6860
rect 10652 6820 15844 6848
rect 10652 6808 10658 6820
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 4246 6780 4252 6792
rect 2898 6752 4252 6780
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 6086 6780 6092 6792
rect 5684 6752 5729 6780
rect 6047 6752 6092 6780
rect 5684 6740 5690 6752
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 6454 6780 6460 6792
rect 6415 6752 6460 6780
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6780 7987 6783
rect 8018 6780 8024 6792
rect 7975 6752 8024 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 8352 6752 9321 6780
rect 8352 6740 8358 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 5353 6715 5411 6721
rect 5353 6681 5365 6715
rect 5399 6712 5411 6715
rect 5399 6684 5580 6712
rect 5399 6681 5411 6684
rect 5353 6675 5411 6681
rect 5552 6656 5580 6684
rect 7190 6672 7196 6724
rect 7248 6672 7254 6724
rect 8938 6712 8944 6724
rect 8899 6684 8944 6712
rect 8938 6672 8944 6684
rect 8996 6672 9002 6724
rect 9122 6712 9128 6724
rect 9083 6684 9128 6712
rect 9122 6672 9128 6684
rect 9180 6672 9186 6724
rect 13262 6672 13268 6724
rect 13320 6712 13326 6724
rect 16114 6712 16120 6724
rect 13320 6684 16120 6712
rect 13320 6672 13326 6684
rect 16114 6672 16120 6684
rect 16172 6672 16178 6724
rect 5534 6604 5540 6656
rect 5592 6604 5598 6656
rect 8389 6647 8447 6653
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 9030 6644 9036 6656
rect 8435 6616 9036 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 15838 6604 15844 6656
rect 15896 6644 15902 6656
rect 16206 6644 16212 6656
rect 15896 6616 16212 6644
rect 15896 6604 15902 6616
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 920 6554 9844 6576
rect 920 6502 3566 6554
rect 3618 6502 3630 6554
rect 3682 6502 3694 6554
rect 3746 6502 3758 6554
rect 3810 6502 3822 6554
rect 3874 6502 8566 6554
rect 8618 6502 8630 6554
rect 8682 6502 8694 6554
rect 8746 6502 8758 6554
rect 8810 6502 8822 6554
rect 8874 6502 9844 6554
rect 920 6480 9844 6502
rect 15470 6468 15476 6520
rect 15528 6508 15534 6520
rect 16206 6508 16212 6520
rect 15528 6480 16212 6508
rect 15528 6468 15534 6480
rect 16206 6468 16212 6480
rect 16264 6468 16270 6520
rect 2222 6440 2228 6452
rect 2183 6412 2228 6440
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 3234 6400 3240 6452
rect 3292 6440 3298 6452
rect 3329 6443 3387 6449
rect 3329 6440 3341 6443
rect 3292 6412 3341 6440
rect 3292 6400 3298 6412
rect 3329 6409 3341 6412
rect 3375 6409 3387 6443
rect 3329 6403 3387 6409
rect 5721 6443 5779 6449
rect 5721 6409 5733 6443
rect 5767 6440 5779 6443
rect 5810 6440 5816 6452
rect 5767 6412 5816 6440
rect 5767 6409 5779 6412
rect 5721 6403 5779 6409
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 7282 6440 7288 6452
rect 6656 6412 7288 6440
rect 4246 6332 4252 6384
rect 4304 6332 4310 6384
rect 4801 6375 4859 6381
rect 4801 6341 4813 6375
rect 4847 6372 4859 6375
rect 5350 6372 5356 6384
rect 4847 6344 5356 6372
rect 4847 6341 4859 6344
rect 4801 6335 4859 6341
rect 5350 6332 5356 6344
rect 5408 6332 5414 6384
rect 6656 6372 6684 6412
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 9122 6440 9128 6452
rect 7524 6412 9128 6440
rect 7524 6400 7530 6412
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 5736 6344 6684 6372
rect 1670 6304 1676 6316
rect 1631 6276 1676 6304
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2409 6307 2467 6313
rect 2409 6304 2421 6307
rect 2188 6276 2421 6304
rect 2188 6264 2194 6276
rect 2409 6273 2421 6276
rect 2455 6273 2467 6307
rect 2409 6267 2467 6273
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 5736 6304 5764 6344
rect 7374 6332 7380 6384
rect 7432 6332 7438 6384
rect 7006 6304 7012 6316
rect 5583 6276 5764 6304
rect 6967 6276 7012 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 5077 6239 5135 6245
rect 5077 6236 5089 6239
rect 5000 6208 5089 6236
rect 1486 6168 1492 6180
rect 1447 6140 1492 6168
rect 1486 6128 1492 6140
rect 1544 6128 1550 6180
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 5000 6100 5028 6208
rect 5077 6205 5089 6208
rect 5123 6236 5135 6239
rect 5626 6236 5632 6248
rect 5123 6208 5632 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 5736 6168 5764 6276
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 8478 6304 8484 6316
rect 8439 6276 8484 6304
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 13872 6276 13952 6304
rect 13872 6264 13878 6276
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6236 6699 6239
rect 6914 6236 6920 6248
rect 6687 6208 6920 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 5644 6140 5764 6168
rect 5644 6112 5672 6140
rect 13924 6112 13952 6276
rect 4120 6072 5028 6100
rect 4120 6060 4126 6072
rect 5626 6060 5632 6112
rect 5684 6060 5690 6112
rect 8938 6100 8944 6112
rect 8899 6072 8944 6100
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 13906 6060 13912 6112
rect 13964 6060 13970 6112
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 7566 6010
rect 7618 5958 7630 6010
rect 7682 5958 7694 6010
rect 7746 5958 7758 6010
rect 7810 5958 7822 6010
rect 7874 5958 9844 6010
rect 13814 5992 13820 6044
rect 13872 6032 13878 6044
rect 14366 6032 14372 6044
rect 13872 6004 14372 6032
rect 13872 5992 13878 6004
rect 14366 5992 14372 6004
rect 14424 5992 14430 6044
rect 16666 5992 16672 6044
rect 16724 5992 16730 6044
rect 920 5936 9844 5958
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 2958 5896 2964 5908
rect 2915 5868 2964 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 5534 5896 5540 5908
rect 5495 5868 5540 5896
rect 5534 5856 5540 5868
rect 5592 5896 5598 5908
rect 6178 5896 6184 5908
rect 5592 5868 6184 5896
rect 5592 5856 5598 5868
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 9122 5896 9128 5908
rect 9083 5868 9128 5896
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 1489 5831 1547 5837
rect 1489 5797 1501 5831
rect 1535 5828 1547 5831
rect 3142 5828 3148 5840
rect 1535 5800 3148 5828
rect 1535 5797 1547 5800
rect 1489 5791 1547 5797
rect 3142 5788 3148 5800
rect 3200 5788 3206 5840
rect 750 5720 756 5772
rect 808 5760 814 5772
rect 808 5732 2176 5760
rect 808 5720 814 5732
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 2038 5692 2044 5704
rect 1443 5664 2044 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2148 5701 2176 5732
rect 2222 5720 2228 5772
rect 2280 5760 2286 5772
rect 3789 5763 3847 5769
rect 2280 5732 2325 5760
rect 2280 5720 2286 5732
rect 3789 5729 3801 5763
rect 3835 5760 3847 5763
rect 4062 5760 4068 5772
rect 3835 5732 4068 5760
rect 3835 5729 3847 5732
rect 3789 5723 3847 5729
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 6822 5760 6828 5772
rect 6783 5732 6828 5760
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 8202 5760 8208 5772
rect 8163 5732 8208 5760
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2774 5692 2780 5704
rect 2363 5664 2780 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3510 5692 3516 5704
rect 3007 5664 3516 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 2056 5624 2084 5652
rect 2682 5624 2688 5636
rect 2056 5596 2688 5624
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 3326 5584 3332 5636
rect 3384 5624 3390 5636
rect 4065 5627 4123 5633
rect 4065 5624 4077 5627
rect 3384 5596 4077 5624
rect 3384 5584 3390 5596
rect 4065 5593 4077 5596
rect 4111 5593 4123 5627
rect 4065 5587 4123 5593
rect 4338 5584 4344 5636
rect 4396 5624 4402 5636
rect 8128 5624 8156 5655
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8444 5664 8953 5692
rect 8444 5652 8450 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 8202 5624 8208 5636
rect 4396 5596 4554 5624
rect 8128 5596 8208 5624
rect 4396 5584 4402 5596
rect 4448 5556 4476 5596
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 16684 5568 16712 5992
rect 5534 5556 5540 5568
rect 4448 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 6822 5516 6828 5568
rect 6880 5556 6886 5568
rect 7374 5556 7380 5568
rect 6880 5528 7380 5556
rect 6880 5516 6886 5528
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 15746 5516 15752 5568
rect 15804 5556 15810 5568
rect 15804 5528 16620 5556
rect 15804 5516 15810 5528
rect 920 5466 9844 5488
rect 920 5414 3566 5466
rect 3618 5414 3630 5466
rect 3682 5414 3694 5466
rect 3746 5414 3758 5466
rect 3810 5414 3822 5466
rect 3874 5414 8566 5466
rect 8618 5414 8630 5466
rect 8682 5414 8694 5466
rect 8746 5414 8758 5466
rect 8810 5414 8822 5466
rect 8874 5414 9844 5466
rect 13538 5448 13544 5500
rect 13596 5488 13602 5500
rect 14182 5488 14188 5500
rect 13596 5460 14188 5488
rect 13596 5448 13602 5460
rect 14182 5448 14188 5460
rect 14240 5448 14246 5500
rect 920 5392 9844 5414
rect 3881 5355 3939 5361
rect 3881 5321 3893 5355
rect 3927 5352 3939 5355
rect 4062 5352 4068 5364
rect 3927 5324 4068 5352
rect 3927 5321 3939 5324
rect 3881 5315 3939 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4617 5355 4675 5361
rect 4617 5321 4629 5355
rect 4663 5352 4675 5355
rect 4890 5352 4896 5364
rect 4663 5324 4896 5352
rect 4663 5321 4675 5324
rect 4617 5315 4675 5321
rect 4890 5312 4896 5324
rect 4948 5312 4954 5364
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 6454 5352 6460 5364
rect 5767 5324 6460 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 6730 5312 6736 5364
rect 6788 5352 6794 5364
rect 6825 5355 6883 5361
rect 6825 5352 6837 5355
rect 6788 5324 6837 5352
rect 6788 5312 6794 5324
rect 6825 5321 6837 5324
rect 6871 5321 6883 5355
rect 6825 5315 6883 5321
rect 566 5244 572 5296
rect 624 5284 630 5296
rect 5810 5284 5816 5296
rect 624 5256 4016 5284
rect 624 5244 630 5256
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 3988 5225 4016 5256
rect 4448 5256 5816 5284
rect 4448 5225 4476 5256
rect 5810 5244 5816 5256
rect 5868 5244 5874 5296
rect 7282 5284 7288 5296
rect 7243 5256 7288 5284
rect 7282 5244 7288 5256
rect 7340 5244 7346 5296
rect 7374 5244 7380 5296
rect 7432 5284 7438 5296
rect 9217 5287 9275 5293
rect 9217 5284 9229 5287
rect 7432 5256 9229 5284
rect 7432 5244 7438 5256
rect 9217 5253 9229 5256
rect 9263 5284 9275 5287
rect 9306 5284 9312 5296
rect 9263 5256 9312 5284
rect 9263 5253 9275 5256
rect 9217 5247 9275 5253
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 2832 5188 3801 5216
rect 2832 5176 2838 5188
rect 3789 5185 3801 5188
rect 3835 5216 3847 5219
rect 3973 5219 4031 5225
rect 3835 5188 3924 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 3896 5080 3924 5188
rect 3973 5185 3985 5219
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 4798 5216 4804 5228
rect 4663 5188 4804 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 6178 5216 6184 5228
rect 6139 5188 6184 5216
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 7300 5216 7328 5244
rect 6788 5188 7328 5216
rect 6788 5176 6794 5188
rect 7466 5176 7472 5228
rect 7524 5216 7530 5228
rect 7524 5188 7617 5216
rect 7524 5176 7530 5188
rect 8570 5176 8576 5228
rect 8628 5216 8634 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8628 5188 8953 5216
rect 8628 5176 8634 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 9030 5176 9036 5228
rect 9088 5216 9094 5228
rect 9088 5188 9133 5216
rect 9088 5176 9094 5188
rect 4154 5108 4160 5160
rect 4212 5148 4218 5160
rect 5077 5151 5135 5157
rect 5077 5148 5089 5151
rect 4212 5120 5089 5148
rect 4212 5108 4218 5120
rect 5077 5117 5089 5120
rect 5123 5117 5135 5151
rect 5077 5111 5135 5117
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 7006 5148 7012 5160
rect 5592 5120 7012 5148
rect 5592 5108 5598 5120
rect 7006 5108 7012 5120
rect 7064 5148 7070 5160
rect 7484 5148 7512 5176
rect 7064 5120 7512 5148
rect 7064 5108 7070 5120
rect 4522 5080 4528 5092
rect 3896 5052 4528 5080
rect 4522 5040 4528 5052
rect 4580 5080 4586 5092
rect 4982 5080 4988 5092
rect 4580 5052 4988 5080
rect 4580 5040 4586 5052
rect 4982 5040 4988 5052
rect 5040 5040 5046 5092
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 7653 5015 7711 5021
rect 7653 5012 7665 5015
rect 7524 4984 7665 5012
rect 7524 4972 7530 4984
rect 7653 4981 7665 4984
rect 7699 4981 7711 5015
rect 7653 4975 7711 4981
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 8941 5015 8999 5021
rect 8941 5012 8953 5015
rect 8352 4984 8953 5012
rect 8352 4972 8358 4984
rect 8941 4981 8953 4984
rect 8987 4981 8999 5015
rect 8941 4975 8999 4981
rect 3036 4922 9844 4944
rect 106 4836 112 4888
rect 164 4876 170 4888
rect 2774 4876 2780 4888
rect 164 4848 2780 4876
rect 164 4836 170 4848
rect 2774 4836 2780 4848
rect 2832 4836 2838 4888
rect 3036 4870 7566 4922
rect 7618 4870 7630 4922
rect 7682 4870 7694 4922
rect 7746 4870 7758 4922
rect 7810 4870 7822 4922
rect 7874 4870 9844 4922
rect 3036 4848 9844 4870
rect 1118 4768 1124 4820
rect 1176 4808 1182 4820
rect 2406 4808 2412 4820
rect 1176 4780 2412 4808
rect 1176 4768 1182 4780
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5997 4811 6055 4817
rect 5997 4808 6009 4811
rect 5592 4780 6009 4808
rect 5592 4768 5598 4780
rect 5997 4777 6009 4780
rect 6043 4777 6055 4811
rect 5997 4771 6055 4777
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 6733 4811 6791 4817
rect 6733 4808 6745 4811
rect 6144 4780 6745 4808
rect 6144 4768 6150 4780
rect 6733 4777 6745 4780
rect 6779 4777 6791 4811
rect 6733 4771 6791 4777
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 6972 4780 7389 4808
rect 6972 4768 6978 4780
rect 7377 4777 7389 4780
rect 7423 4777 7435 4811
rect 8386 4808 8392 4820
rect 8347 4780 8392 4808
rect 7377 4771 7435 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 934 4700 940 4752
rect 992 4740 998 4752
rect 4154 4740 4160 4752
rect 992 4712 4160 4740
rect 992 4700 998 4712
rect 4154 4700 4160 4712
rect 4212 4700 4218 4752
rect 1118 4632 1124 4684
rect 1176 4672 1182 4684
rect 1302 4672 1308 4684
rect 1176 4644 1308 4672
rect 1176 4632 1182 4644
rect 1302 4632 1308 4644
rect 1360 4632 1366 4684
rect 3418 4632 3424 4684
rect 3476 4672 3482 4684
rect 4890 4672 4896 4684
rect 3476 4644 4384 4672
rect 4851 4644 4896 4672
rect 3476 4632 3482 4644
rect 1210 4564 1216 4616
rect 1268 4564 1274 4616
rect 1854 4564 1860 4616
rect 1912 4604 1918 4616
rect 2866 4604 2872 4616
rect 1912 4576 2872 4604
rect 1912 4564 1918 4576
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3694 4604 3700 4616
rect 3655 4576 3700 4604
rect 3513 4567 3571 4573
rect 1228 4536 1256 4564
rect 3528 4536 3556 4567
rect 3694 4564 3700 4576
rect 3752 4564 3758 4616
rect 4356 4613 4384 4644
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 6638 4672 6644 4684
rect 6196 4644 6644 4672
rect 6196 4613 6224 4644
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 8386 4632 8392 4684
rect 8444 4672 8450 4684
rect 9306 4672 9312 4684
rect 8444 4644 9312 4672
rect 8444 4632 8450 4644
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6270 4564 6276 4616
rect 6328 4604 6334 4616
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 6328 4576 6837 4604
rect 6328 4564 6334 4576
rect 6825 4573 6837 4576
rect 6871 4604 6883 4607
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 6871 4576 7297 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 7285 4573 7297 4576
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 8938 4604 8944 4616
rect 8619 4576 8944 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 9232 4613 9260 4644
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 4062 4536 4068 4548
rect 1228 4508 2774 4536
rect 3528 4508 4068 4536
rect 2746 4128 2774 4508
rect 4062 4496 4068 4508
rect 4120 4496 4126 4548
rect 9306 4536 9312 4548
rect 9267 4508 9312 4536
rect 9306 4496 9312 4508
rect 9364 4496 9370 4548
rect 3697 4471 3755 4477
rect 3697 4437 3709 4471
rect 3743 4468 3755 4471
rect 4246 4468 4252 4480
rect 3743 4440 4252 4468
rect 3743 4437 3755 4440
rect 3697 4431 3755 4437
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 3036 4378 9844 4400
rect 3036 4326 3566 4378
rect 3618 4326 3630 4378
rect 3682 4326 3694 4378
rect 3746 4326 3758 4378
rect 3810 4326 3822 4378
rect 3874 4326 8566 4378
rect 8618 4326 8630 4378
rect 8682 4326 8694 4378
rect 8746 4326 8758 4378
rect 8810 4326 8822 4378
rect 8874 4326 9844 4378
rect 3036 4304 9844 4326
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 4893 4267 4951 4273
rect 4893 4264 4905 4267
rect 4488 4236 4905 4264
rect 4488 4224 4494 4236
rect 4893 4233 4905 4236
rect 4939 4233 4951 4267
rect 4893 4227 4951 4233
rect 8202 4224 8208 4276
rect 8260 4224 8266 4276
rect 8220 4196 8248 4224
rect 6840 4168 8248 4196
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 2746 4100 3709 4128
rect 3697 4097 3709 4100
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4890 4128 4896 4140
rect 4212 4100 4896 4128
rect 4212 4088 4218 4100
rect 4890 4088 4896 4100
rect 4948 4128 4954 4140
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4948 4100 4997 4128
rect 4948 4088 4954 4100
rect 4985 4097 4997 4100
rect 5031 4128 5043 4131
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 5031 4100 5457 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 5445 4091 5503 4097
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4128 6147 4131
rect 6840 4128 6868 4168
rect 6135 4100 6868 4128
rect 6917 4131 6975 4137
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 6917 4097 6929 4131
rect 6963 4128 6975 4131
rect 7006 4128 7012 4140
rect 6963 4100 7012 4128
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4128 7895 4131
rect 8202 4128 8208 4140
rect 7883 4100 8208 4128
rect 7883 4097 7895 4100
rect 7837 4091 7895 4097
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4128 9091 4131
rect 9214 4128 9220 4140
rect 9079 4100 9220 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 12434 4128 12440 4140
rect 12400 4100 12440 4128
rect 12400 4088 12406 4100
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 4062 4060 4068 4072
rect 4023 4032 4068 4060
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 6546 4020 6552 4072
rect 6604 4060 6610 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6604 4032 6837 4060
rect 6604 4020 6610 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 6270 3992 6276 4004
rect 6231 3964 6276 3992
rect 6270 3952 6276 3964
rect 6328 3952 6334 4004
rect 5534 3924 5540 3936
rect 5495 3896 5540 3924
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 7340 3896 7757 3924
rect 7340 3884 7346 3896
rect 7745 3893 7757 3896
rect 7791 3893 7803 3927
rect 9214 3924 9220 3936
rect 9175 3896 9220 3924
rect 7745 3887 7803 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 3036 3834 9844 3856
rect 3036 3782 7566 3834
rect 7618 3782 7630 3834
rect 7682 3782 7694 3834
rect 7746 3782 7758 3834
rect 7810 3782 7822 3834
rect 7874 3782 9844 3834
rect 3036 3760 9844 3782
rect 3697 3723 3755 3729
rect 3697 3689 3709 3723
rect 3743 3689 3755 3723
rect 3697 3683 3755 3689
rect 4249 3723 4307 3729
rect 4249 3689 4261 3723
rect 4295 3720 4307 3723
rect 4614 3720 4620 3732
rect 4295 3692 4620 3720
rect 4295 3689 4307 3692
rect 4249 3683 4307 3689
rect 3712 3652 3740 3683
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 4893 3723 4951 3729
rect 4893 3689 4905 3723
rect 4939 3720 4951 3723
rect 5074 3720 5080 3732
rect 4939 3692 5080 3720
rect 4939 3689 4951 3692
rect 4893 3683 4951 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 6086 3720 6092 3732
rect 6047 3692 6092 3720
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 6822 3720 6828 3732
rect 6783 3692 6828 3720
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7190 3680 7196 3732
rect 7248 3720 7254 3732
rect 7469 3723 7527 3729
rect 7469 3720 7481 3723
rect 7248 3692 7481 3720
rect 7248 3680 7254 3692
rect 7469 3689 7481 3692
rect 7515 3689 7527 3723
rect 8018 3720 8024 3732
rect 7979 3692 8024 3720
rect 7469 3683 7527 3689
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 5166 3652 5172 3664
rect 3712 3624 5172 3652
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 9398 3584 9404 3596
rect 6604 3556 6960 3584
rect 6604 3544 6610 3556
rect 3510 3516 3516 3528
rect 3471 3488 3516 3516
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 4154 3516 4160 3528
rect 4115 3488 4160 3516
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4522 3516 4528 3528
rect 4387 3488 4528 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 4706 3476 4712 3528
rect 4764 3516 4770 3528
rect 4801 3519 4859 3525
rect 4801 3516 4813 3519
rect 4764 3488 4813 3516
rect 4764 3476 4770 3488
rect 4801 3485 4813 3488
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3485 5043 3519
rect 5902 3516 5908 3528
rect 5863 3488 5908 3516
rect 4985 3479 5043 3485
rect 4540 3448 4568 3476
rect 5000 3448 5028 3479
rect 5902 3476 5908 3488
rect 5960 3476 5966 3528
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 6932 3525 6960 3556
rect 8220 3556 9404 3584
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6696 3488 6745 3516
rect 6696 3476 6702 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 6917 3519 6975 3525
rect 6917 3485 6929 3519
rect 6963 3516 6975 3519
rect 7377 3519 7435 3525
rect 7377 3516 7389 3519
rect 6963 3488 7389 3516
rect 6963 3485 6975 3488
rect 6917 3479 6975 3485
rect 7377 3485 7389 3488
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3516 7619 3519
rect 8110 3516 8116 3528
rect 7607 3488 8116 3516
rect 7607 3485 7619 3488
rect 7561 3479 7619 3485
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 8220 3525 8248 3556
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 9033 3519 9091 3525
rect 9033 3485 9045 3519
rect 9079 3516 9091 3519
rect 9122 3516 9128 3528
rect 9079 3488 9128 3516
rect 9079 3485 9091 3488
rect 9033 3479 9091 3485
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 5074 3448 5080 3460
rect 4540 3420 5080 3448
rect 5074 3408 5080 3420
rect 5132 3448 5138 3460
rect 5718 3448 5724 3460
rect 5132 3420 5724 3448
rect 5132 3408 5138 3420
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 10318 3408 10324 3460
rect 10376 3448 10382 3460
rect 16206 3448 16212 3460
rect 10376 3420 16212 3448
rect 10376 3408 10382 3420
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 9214 3380 9220 3392
rect 9175 3352 9220 3380
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 3036 3290 9844 3312
rect 3036 3238 3566 3290
rect 3618 3238 3630 3290
rect 3682 3238 3694 3290
rect 3746 3238 3758 3290
rect 3810 3238 3822 3290
rect 3874 3238 8566 3290
rect 8618 3238 8630 3290
rect 8682 3238 8694 3290
rect 8746 3238 8758 3290
rect 8810 3238 8822 3290
rect 8874 3238 9844 3290
rect 3036 3216 9844 3238
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 3697 3179 3755 3185
rect 3697 3176 3709 3179
rect 3292 3148 3709 3176
rect 3292 3136 3298 3148
rect 3697 3145 3709 3148
rect 3743 3145 3755 3179
rect 4982 3176 4988 3188
rect 4943 3148 4988 3176
rect 3697 3139 3755 3145
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 5721 3179 5779 3185
rect 5721 3145 5733 3179
rect 5767 3176 5779 3179
rect 5994 3176 6000 3188
rect 5767 3148 6000 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6181 3179 6239 3185
rect 6181 3145 6193 3179
rect 6227 3176 6239 3179
rect 6730 3176 6736 3188
rect 6227 3148 6736 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 6914 3176 6920 3188
rect 6875 3148 6920 3176
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 7929 3179 7987 3185
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 8478 3176 8484 3188
rect 7975 3148 8484 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 9214 3176 9220 3188
rect 9175 3148 9220 3176
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 5626 3108 5632 3120
rect 4356 3080 5632 3108
rect 3510 3040 3516 3052
rect 3471 3012 3516 3040
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3040 4215 3043
rect 4246 3040 4252 3052
rect 4203 3012 4252 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4356 3049 4384 3080
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 13906 3108 13912 3120
rect 6380 3080 13912 3108
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 4890 3040 4896 3052
rect 4488 3012 4896 3040
rect 4488 3000 4494 3012
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 5534 3040 5540 3052
rect 5495 3012 5540 3040
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 5718 3040 5724 3052
rect 5679 3012 5724 3040
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 6380 3049 6408 3080
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 4908 2972 4936 3000
rect 6840 2972 6868 3003
rect 7466 3000 7472 3052
rect 7524 3040 7530 3052
rect 7745 3043 7803 3049
rect 7745 3040 7757 3043
rect 7524 3012 7757 3040
rect 7524 3000 7530 3012
rect 7745 3009 7757 3012
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9766 3040 9772 3052
rect 9079 3012 9772 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9766 3000 9772 3012
rect 9824 3000 9830 3052
rect 4908 2944 6868 2972
rect 14090 2864 14096 2916
rect 14148 2904 14154 2916
rect 16390 2904 16396 2916
rect 14148 2876 16396 2904
rect 14148 2864 14154 2876
rect 16390 2864 16396 2876
rect 16448 2864 16454 2916
rect 3878 2796 3884 2848
rect 3936 2836 3942 2848
rect 4157 2839 4215 2845
rect 4157 2836 4169 2839
rect 3936 2808 4169 2836
rect 3936 2796 3942 2808
rect 4157 2805 4169 2808
rect 4203 2805 4215 2839
rect 4157 2799 4215 2805
rect 3036 2746 9844 2768
rect 3036 2694 7566 2746
rect 7618 2694 7630 2746
rect 7682 2694 7694 2746
rect 7746 2694 7758 2746
rect 7810 2694 7822 2746
rect 7874 2694 9844 2746
rect 3036 2672 9844 2694
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4249 2635 4307 2641
rect 4249 2632 4261 2635
rect 4212 2604 4261 2632
rect 4212 2592 4218 2604
rect 4249 2601 4261 2604
rect 4295 2601 4307 2635
rect 4249 2595 4307 2601
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 8018 2632 8024 2644
rect 6595 2604 8024 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 9030 2632 9036 2644
rect 8527 2604 9036 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 2774 2456 2780 2508
rect 2832 2456 2838 2508
rect 7374 2496 7380 2508
rect 5920 2468 7380 2496
rect 2792 2428 2820 2456
rect 3697 2431 3755 2437
rect 3697 2428 3709 2431
rect 2792 2400 3709 2428
rect 3697 2397 3709 2400
rect 3743 2428 3755 2431
rect 4157 2431 4215 2437
rect 4157 2428 4169 2431
rect 3743 2400 4169 2428
rect 3743 2397 3755 2400
rect 3697 2391 3755 2397
rect 4157 2397 4169 2400
rect 4203 2397 4215 2431
rect 4157 2391 4215 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4580 2400 4813 2428
rect 4580 2388 4586 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5074 2428 5080 2440
rect 5031 2400 5080 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5074 2388 5080 2400
rect 5132 2388 5138 2440
rect 5920 2437 5948 2468
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 9398 2496 9404 2508
rect 8404 2468 9404 2496
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 6730 2428 6736 2440
rect 6691 2400 6736 2428
rect 5905 2391 5963 2397
rect 6730 2388 6736 2400
rect 6788 2388 6794 2440
rect 8404 2437 8432 2468
rect 9398 2456 9404 2468
rect 9456 2456 9462 2508
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 8536 2400 8585 2428
rect 8536 2388 8542 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 9950 2428 9956 2440
rect 9263 2400 9956 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 3142 2252 3148 2304
rect 3200 2292 3206 2304
rect 3605 2295 3663 2301
rect 3605 2292 3617 2295
rect 3200 2264 3617 2292
rect 3200 2252 3206 2264
rect 3605 2261 3617 2264
rect 3651 2261 3663 2295
rect 4890 2292 4896 2304
rect 4851 2264 4896 2292
rect 3605 2255 3663 2261
rect 4890 2252 4896 2264
rect 4948 2252 4954 2304
rect 5994 2292 6000 2304
rect 5955 2264 6000 2292
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 8110 2252 8116 2304
rect 8168 2292 8174 2304
rect 9033 2295 9091 2301
rect 9033 2292 9045 2295
rect 8168 2264 9045 2292
rect 8168 2252 8174 2264
rect 9033 2261 9045 2264
rect 9079 2261 9091 2295
rect 9033 2255 9091 2261
rect 3036 2202 9844 2224
rect 3036 2150 3566 2202
rect 3618 2150 3630 2202
rect 3682 2150 3694 2202
rect 3746 2150 3758 2202
rect 3810 2150 3822 2202
rect 3874 2150 8566 2202
rect 8618 2150 8630 2202
rect 8682 2150 8694 2202
rect 8746 2150 8758 2202
rect 8810 2150 8822 2202
rect 8874 2150 9844 2202
rect 3036 2128 9844 2150
rect 3326 2048 3332 2100
rect 3384 2088 3390 2100
rect 3605 2091 3663 2097
rect 3605 2088 3617 2091
rect 3384 2060 3617 2088
rect 3384 2048 3390 2060
rect 3605 2057 3617 2060
rect 3651 2057 3663 2091
rect 5442 2088 5448 2100
rect 3605 2051 3663 2057
rect 4172 2060 5448 2088
rect 4062 2020 4068 2032
rect 3528 1992 4068 2020
rect 3528 1961 3556 1992
rect 4062 1980 4068 1992
rect 4120 1980 4126 2032
rect 3513 1955 3571 1961
rect 3513 1921 3525 1955
rect 3559 1921 3571 1955
rect 3513 1915 3571 1921
rect 3697 1955 3755 1961
rect 3697 1921 3709 1955
rect 3743 1952 3755 1955
rect 3970 1952 3976 1964
rect 3743 1924 3976 1952
rect 3743 1921 3755 1924
rect 3697 1915 3755 1921
rect 3970 1912 3976 1924
rect 4028 1912 4034 1964
rect 4172 1961 4200 2060
rect 5442 2048 5448 2060
rect 5500 2048 5506 2100
rect 5626 2088 5632 2100
rect 5587 2060 5632 2088
rect 5626 2048 5632 2060
rect 5684 2048 5690 2100
rect 8478 2048 8484 2100
rect 8536 2088 8542 2100
rect 8573 2091 8631 2097
rect 8573 2088 8585 2091
rect 8536 2060 8585 2088
rect 8536 2048 8542 2060
rect 8573 2057 8585 2060
rect 8619 2057 8631 2091
rect 8573 2051 8631 2057
rect 9217 2091 9275 2097
rect 9217 2057 9229 2091
rect 9263 2088 9275 2091
rect 9490 2088 9496 2100
rect 9263 2060 9496 2088
rect 9263 2057 9275 2060
rect 9217 2051 9275 2057
rect 9490 2048 9496 2060
rect 9548 2048 9554 2100
rect 4338 1980 4344 2032
rect 4396 2020 4402 2032
rect 4893 2023 4951 2029
rect 4893 2020 4905 2023
rect 4396 1992 4905 2020
rect 4396 1980 4402 1992
rect 4893 1989 4905 1992
rect 4939 1989 4951 2023
rect 4893 1983 4951 1989
rect 5994 1980 6000 2032
rect 6052 2020 6058 2032
rect 9030 2020 9036 2032
rect 6052 1992 9036 2020
rect 6052 1980 6058 1992
rect 4157 1955 4215 1961
rect 4157 1921 4169 1955
rect 4203 1921 4215 1955
rect 4798 1952 4804 1964
rect 4759 1924 4804 1952
rect 4157 1915 4215 1921
rect 4798 1912 4804 1924
rect 4856 1912 4862 1964
rect 4985 1955 5043 1961
rect 4985 1921 4997 1955
rect 5031 1952 5043 1955
rect 5074 1952 5080 1964
rect 5031 1924 5080 1952
rect 5031 1921 5043 1924
rect 4985 1915 5043 1921
rect 5074 1912 5080 1924
rect 5132 1912 5138 1964
rect 5442 1952 5448 1964
rect 5403 1924 5448 1952
rect 5442 1912 5448 1924
rect 5500 1912 5506 1964
rect 5629 1955 5687 1961
rect 5629 1921 5641 1955
rect 5675 1921 5687 1955
rect 6086 1952 6092 1964
rect 6047 1924 6092 1952
rect 5629 1915 5687 1921
rect 5092 1884 5120 1912
rect 5644 1884 5672 1915
rect 6086 1912 6092 1924
rect 6144 1912 6150 1964
rect 6748 1961 6776 1992
rect 9030 1980 9036 1992
rect 9088 1980 9094 2032
rect 6733 1955 6791 1961
rect 6733 1921 6745 1955
rect 6779 1921 6791 1955
rect 6914 1952 6920 1964
rect 6875 1924 6920 1952
rect 6733 1915 6791 1921
rect 6914 1912 6920 1924
rect 6972 1912 6978 1964
rect 8665 1955 8723 1961
rect 8665 1921 8677 1955
rect 8711 1952 8723 1955
rect 9214 1952 9220 1964
rect 8711 1924 9220 1952
rect 8711 1921 8723 1924
rect 8665 1915 8723 1921
rect 9214 1912 9220 1924
rect 9272 1912 9278 1964
rect 9309 1955 9367 1961
rect 9309 1921 9321 1955
rect 9355 1952 9367 1955
rect 9582 1952 9588 1964
rect 9355 1924 9588 1952
rect 9355 1921 9367 1924
rect 9309 1915 9367 1921
rect 9582 1912 9588 1924
rect 9640 1912 9646 1964
rect 5092 1856 5672 1884
rect 4246 1816 4252 1828
rect 4207 1788 4252 1816
rect 4246 1776 4252 1788
rect 4304 1776 4310 1828
rect 6270 1748 6276 1760
rect 6231 1720 6276 1748
rect 6270 1708 6276 1720
rect 6328 1708 6334 1760
rect 6822 1748 6828 1760
rect 6783 1720 6828 1748
rect 6822 1708 6828 1720
rect 6880 1708 6886 1760
rect 3036 1658 9844 1680
rect 3036 1606 7566 1658
rect 7618 1606 7630 1658
rect 7682 1606 7694 1658
rect 7746 1606 7758 1658
rect 7810 1606 7822 1658
rect 7874 1606 9844 1658
rect 3036 1584 9844 1606
rect 16592 1612 16620 5528
rect 16666 5516 16672 5568
rect 16724 5516 16730 5568
rect 16666 1612 16672 1624
rect 16592 1584 16672 1612
rect 16666 1572 16672 1584
rect 16724 1572 16730 1624
rect 658 1504 664 1556
rect 716 1544 722 1556
rect 4890 1544 4896 1556
rect 716 1516 4896 1544
rect 716 1504 722 1516
rect 4890 1504 4896 1516
rect 4948 1504 4954 1556
rect 198 1436 204 1488
rect 256 1476 262 1488
rect 4798 1476 4804 1488
rect 256 1448 4804 1476
rect 256 1436 262 1448
rect 4798 1436 4804 1448
rect 4856 1436 4862 1488
rect 8938 1476 8944 1488
rect 8899 1448 8944 1476
rect 8938 1436 8944 1448
rect 8996 1436 9002 1488
rect 382 1368 388 1420
rect 440 1408 446 1420
rect 5442 1408 5448 1420
rect 440 1380 5448 1408
rect 440 1368 446 1380
rect 5442 1368 5448 1380
rect 5500 1368 5506 1420
rect 6822 1368 6828 1420
rect 6880 1408 6886 1420
rect 6880 1380 6960 1408
rect 6880 1368 6886 1380
rect 2958 1300 2964 1352
rect 3016 1340 3022 1352
rect 3513 1343 3571 1349
rect 3513 1340 3525 1343
rect 3016 1312 3525 1340
rect 3016 1300 3022 1312
rect 3513 1309 3525 1312
rect 3559 1309 3571 1343
rect 3513 1303 3571 1309
rect 4341 1343 4399 1349
rect 4341 1309 4353 1343
rect 4387 1340 4399 1343
rect 4430 1340 4436 1352
rect 4387 1312 4436 1340
rect 4387 1309 4399 1312
rect 4341 1303 4399 1309
rect 4430 1300 4436 1312
rect 4488 1300 4494 1352
rect 4798 1340 4804 1352
rect 4759 1312 4804 1340
rect 4798 1300 4804 1312
rect 4856 1300 4862 1352
rect 4985 1343 5043 1349
rect 4985 1309 4997 1343
rect 5031 1340 5043 1343
rect 5074 1340 5080 1352
rect 5031 1312 5080 1340
rect 5031 1309 5043 1312
rect 4985 1303 5043 1309
rect 5074 1300 5080 1312
rect 5132 1300 5138 1352
rect 5258 1300 5264 1352
rect 5316 1340 5322 1352
rect 5905 1343 5963 1349
rect 5905 1340 5917 1343
rect 5316 1312 5917 1340
rect 5316 1300 5322 1312
rect 5905 1309 5917 1312
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 6089 1343 6147 1349
rect 6089 1309 6101 1343
rect 6135 1309 6147 1343
rect 6730 1340 6736 1352
rect 6691 1312 6736 1340
rect 6089 1303 6147 1309
rect 4246 1272 4252 1284
rect 4207 1244 4252 1272
rect 4246 1232 4252 1244
rect 4304 1232 4310 1284
rect 5092 1272 5120 1300
rect 6104 1272 6132 1303
rect 6730 1300 6736 1312
rect 6788 1300 6794 1352
rect 6932 1340 6960 1380
rect 7193 1343 7251 1349
rect 7193 1340 7205 1343
rect 6932 1312 7205 1340
rect 7193 1309 7205 1312
rect 7239 1309 7251 1343
rect 7193 1303 7251 1309
rect 7377 1343 7435 1349
rect 7377 1309 7389 1343
rect 7423 1340 7435 1343
rect 8202 1340 8208 1352
rect 7423 1312 8208 1340
rect 7423 1309 7435 1312
rect 7377 1303 7435 1309
rect 8202 1300 8208 1312
rect 8260 1300 8266 1352
rect 5092 1244 6132 1272
rect 3697 1207 3755 1213
rect 3697 1173 3709 1207
rect 3743 1204 3755 1207
rect 4062 1204 4068 1216
rect 3743 1176 4068 1204
rect 3743 1173 3755 1176
rect 3697 1167 3755 1173
rect 4062 1164 4068 1176
rect 4120 1164 4126 1216
rect 4982 1204 4988 1216
rect 4943 1176 4988 1204
rect 4982 1164 4988 1176
rect 5040 1164 5046 1216
rect 6086 1204 6092 1216
rect 6047 1176 6092 1204
rect 6086 1164 6092 1176
rect 6144 1164 6150 1216
rect 6546 1204 6552 1216
rect 6507 1176 6552 1204
rect 6546 1164 6552 1176
rect 6604 1164 6610 1216
rect 7374 1204 7380 1216
rect 7335 1176 7380 1204
rect 7374 1164 7380 1176
rect 7432 1164 7438 1216
rect 9122 1204 9128 1216
rect 9083 1176 9128 1204
rect 9122 1164 9128 1176
rect 9180 1164 9186 1216
rect 3036 1114 9844 1136
rect 3036 1062 3566 1114
rect 3618 1062 3630 1114
rect 3682 1062 3694 1114
rect 3746 1062 3758 1114
rect 3810 1062 3822 1114
rect 3874 1062 8566 1114
rect 8618 1062 8630 1114
rect 8682 1062 8694 1114
rect 8746 1062 8758 1114
rect 8810 1062 8822 1114
rect 8874 1062 9844 1114
rect 3036 1040 9844 1062
<< via1 >>
rect 3240 15852 3292 15904
rect 8484 15852 8536 15904
rect 2566 15750 2618 15802
rect 2630 15750 2682 15802
rect 2694 15750 2746 15802
rect 2758 15750 2810 15802
rect 2822 15750 2874 15802
rect 7566 15750 7618 15802
rect 7630 15750 7682 15802
rect 7694 15750 7746 15802
rect 7758 15750 7810 15802
rect 7822 15750 7874 15802
rect 4068 15648 4120 15700
rect 9128 15691 9180 15700
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 8116 15555 8168 15564
rect 8116 15521 8125 15555
rect 8125 15521 8159 15555
rect 8159 15521 8168 15555
rect 8116 15512 8168 15521
rect 2688 15444 2740 15496
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 5724 15487 5776 15496
rect 5724 15453 5733 15487
rect 5733 15453 5767 15487
rect 5767 15453 5776 15487
rect 5724 15444 5776 15453
rect 8392 15487 8444 15496
rect 8392 15453 8401 15487
rect 8401 15453 8435 15487
rect 8435 15453 8444 15487
rect 8392 15444 8444 15453
rect 1400 15376 1452 15428
rect 2136 15376 2188 15428
rect 3148 15376 3200 15428
rect 4620 15419 4672 15428
rect 4620 15385 4629 15419
rect 4629 15385 4663 15419
rect 4663 15385 4672 15419
rect 4620 15376 4672 15385
rect 7380 15376 7432 15428
rect 8024 15376 8076 15428
rect 16672 15376 16724 15428
rect 1216 15308 1268 15360
rect 5540 15308 5592 15360
rect 3566 15206 3618 15258
rect 3630 15206 3682 15258
rect 3694 15206 3746 15258
rect 3758 15206 3810 15258
rect 3822 15206 3874 15258
rect 8566 15206 8618 15258
rect 8630 15206 8682 15258
rect 8694 15206 8746 15258
rect 8758 15206 8810 15258
rect 8822 15206 8874 15258
rect 5724 15104 5776 15156
rect 15384 15104 15436 15156
rect 16580 15104 16632 15156
rect 480 15036 532 15088
rect 4068 15036 4120 15088
rect 7380 15036 7432 15088
rect 8208 15036 8260 15088
rect 3148 14968 3200 15020
rect 9864 14968 9916 15020
rect 16580 14968 16632 15020
rect 2964 14900 3016 14952
rect 4252 14900 4304 14952
rect 4344 14943 4396 14952
rect 4344 14909 4353 14943
rect 4353 14909 4387 14943
rect 4387 14909 4396 14943
rect 5356 14943 5408 14952
rect 4344 14900 4396 14909
rect 5356 14909 5365 14943
rect 5365 14909 5399 14943
rect 5399 14909 5408 14943
rect 5356 14900 5408 14909
rect 8392 14943 8444 14952
rect 8392 14909 8401 14943
rect 8401 14909 8435 14943
rect 8435 14909 8444 14943
rect 8392 14900 8444 14909
rect 296 14832 348 14884
rect 2780 14832 2832 14884
rect 3240 14832 3292 14884
rect 4804 14875 4856 14884
rect 4804 14841 4813 14875
rect 4813 14841 4847 14875
rect 4847 14841 4856 14875
rect 4804 14832 4856 14841
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 3884 14764 3936 14816
rect 9220 14807 9272 14816
rect 9220 14773 9229 14807
rect 9229 14773 9263 14807
rect 9263 14773 9272 14807
rect 9220 14764 9272 14773
rect 2566 14662 2618 14714
rect 2630 14662 2682 14714
rect 2694 14662 2746 14714
rect 2758 14662 2810 14714
rect 2822 14662 2874 14714
rect 7566 14662 7618 14714
rect 7630 14662 7682 14714
rect 7694 14662 7746 14714
rect 7758 14662 7810 14714
rect 7822 14662 7874 14714
rect 756 14560 808 14612
rect 3240 14467 3292 14476
rect 3240 14433 3249 14467
rect 3249 14433 3283 14467
rect 3283 14433 3292 14467
rect 3240 14424 3292 14433
rect 4068 14424 4120 14476
rect 5448 14424 5500 14476
rect 8208 14356 8260 14408
rect 2504 14288 2556 14340
rect 5356 14288 5408 14340
rect 7012 14331 7064 14340
rect 7012 14297 7021 14331
rect 7021 14297 7055 14331
rect 7055 14297 7064 14331
rect 7012 14288 7064 14297
rect 8392 14288 8444 14340
rect 9220 14288 9272 14340
rect 1584 14220 1636 14272
rect 3148 14220 3200 14272
rect 4068 14220 4120 14272
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 7104 14220 7156 14272
rect 9312 14263 9364 14272
rect 9312 14229 9321 14263
rect 9321 14229 9355 14263
rect 9355 14229 9364 14263
rect 9312 14220 9364 14229
rect 3566 14118 3618 14170
rect 3630 14118 3682 14170
rect 3694 14118 3746 14170
rect 3758 14118 3810 14170
rect 3822 14118 3874 14170
rect 8566 14118 8618 14170
rect 8630 14118 8682 14170
rect 8694 14118 8746 14170
rect 8758 14118 8810 14170
rect 8822 14118 8874 14170
rect 3608 14016 3660 14068
rect 4804 14016 4856 14068
rect 5724 14059 5776 14068
rect 5724 14025 5733 14059
rect 5733 14025 5767 14059
rect 5767 14025 5776 14059
rect 5724 14016 5776 14025
rect 3332 13948 3384 14000
rect 5264 13948 5316 14000
rect 9220 14016 9272 14068
rect 8116 13948 8168 14000
rect 1308 13880 1360 13932
rect 4436 13923 4488 13932
rect 4436 13889 4445 13923
rect 4445 13889 4479 13923
rect 4479 13889 4488 13923
rect 4436 13880 4488 13889
rect 6644 13923 6696 13932
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 2044 13812 2096 13864
rect 2412 13812 2464 13864
rect 3608 13812 3660 13864
rect 4896 13855 4948 13864
rect 4896 13821 4905 13855
rect 4905 13821 4939 13855
rect 4939 13821 4948 13855
rect 4896 13812 4948 13821
rect 4712 13744 4764 13796
rect 6644 13889 6653 13923
rect 6653 13889 6687 13923
rect 6687 13889 6696 13923
rect 6644 13880 6696 13889
rect 7104 13880 7156 13932
rect 9588 13880 9640 13932
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 8944 13812 8996 13821
rect 2566 13574 2618 13626
rect 2630 13574 2682 13626
rect 2694 13574 2746 13626
rect 2758 13574 2810 13626
rect 2822 13574 2874 13626
rect 7566 13574 7618 13626
rect 7630 13574 7682 13626
rect 7694 13574 7746 13626
rect 7758 13574 7810 13626
rect 7822 13574 7874 13626
rect 8024 13472 8076 13524
rect 4160 13336 4212 13388
rect 5264 13336 5316 13388
rect 5724 13336 5776 13388
rect 16120 13336 16172 13388
rect 16672 13336 16724 13388
rect 3240 13268 3292 13320
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 7932 13268 7984 13320
rect 8944 13311 8996 13320
rect 2320 13200 2372 13252
rect 6644 13200 6696 13252
rect 6920 13200 6972 13252
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 8944 13268 8996 13277
rect 10140 13268 10192 13320
rect 14280 13268 14332 13320
rect 940 13132 992 13184
rect 8208 13175 8260 13184
rect 8208 13141 8217 13175
rect 8217 13141 8251 13175
rect 8251 13141 8260 13175
rect 8208 13132 8260 13141
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 3566 13030 3618 13082
rect 3630 13030 3682 13082
rect 3694 13030 3746 13082
rect 3758 13030 3810 13082
rect 3822 13030 3874 13082
rect 8566 13030 8618 13082
rect 8630 13030 8682 13082
rect 8694 13030 8746 13082
rect 8758 13030 8810 13082
rect 8822 13030 8874 13082
rect 8300 12971 8352 12980
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 10324 12928 10376 12980
rect 15752 12928 15804 12980
rect 3884 12860 3936 12912
rect 7288 12860 7340 12912
rect 1584 12792 1636 12844
rect 2412 12792 2464 12844
rect 4344 12835 4396 12844
rect 4344 12801 4353 12835
rect 4353 12801 4387 12835
rect 4387 12801 4396 12835
rect 4344 12792 4396 12801
rect 5448 12792 5500 12844
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 2504 12767 2556 12776
rect 2504 12733 2513 12767
rect 2513 12733 2547 12767
rect 2547 12733 2556 12767
rect 2504 12724 2556 12733
rect 5816 12724 5868 12776
rect 6368 12724 6420 12776
rect 7196 12724 7248 12776
rect 9956 12724 10008 12776
rect 16028 12724 16080 12776
rect 112 12588 164 12640
rect 4804 12631 4856 12640
rect 4804 12597 4813 12631
rect 4813 12597 4847 12631
rect 4847 12597 4856 12631
rect 4804 12588 4856 12597
rect 7288 12588 7340 12640
rect 7932 12588 7984 12640
rect 9588 12588 9640 12640
rect 2566 12486 2618 12538
rect 2630 12486 2682 12538
rect 2694 12486 2746 12538
rect 2758 12486 2810 12538
rect 2822 12486 2874 12538
rect 7566 12486 7618 12538
rect 7630 12486 7682 12538
rect 7694 12486 7746 12538
rect 7758 12486 7810 12538
rect 7822 12486 7874 12538
rect 6828 12384 6880 12436
rect 9128 12384 9180 12436
rect 16396 12384 16448 12436
rect 13820 12316 13872 12368
rect 14280 12316 14332 12368
rect 2964 12248 3016 12300
rect 3332 12180 3384 12232
rect 7196 12248 7248 12300
rect 8116 12248 8168 12300
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 4712 12180 4764 12232
rect 6828 12180 6880 12232
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 9036 12180 9088 12232
rect 2688 12112 2740 12164
rect 1584 12044 1636 12096
rect 2044 12044 2096 12096
rect 5724 12112 5776 12164
rect 4068 12044 4120 12096
rect 6920 12044 6972 12096
rect 9772 12044 9824 12096
rect 16212 12044 16264 12096
rect 16396 12044 16448 12096
rect 3566 11942 3618 11994
rect 3630 11942 3682 11994
rect 3694 11942 3746 11994
rect 3758 11942 3810 11994
rect 3822 11942 3874 11994
rect 8566 11942 8618 11994
rect 8630 11942 8682 11994
rect 8694 11942 8746 11994
rect 8758 11942 8810 11994
rect 8822 11942 8874 11994
rect 10508 11908 10560 11960
rect 16212 11908 16264 11960
rect 2688 11772 2740 11824
rect 3332 11772 3384 11824
rect 5816 11815 5868 11824
rect 3332 11679 3384 11688
rect 3332 11645 3341 11679
rect 3341 11645 3375 11679
rect 3375 11645 3384 11679
rect 3332 11636 3384 11645
rect 5816 11781 5825 11815
rect 5825 11781 5859 11815
rect 5859 11781 5868 11815
rect 5816 11772 5868 11781
rect 7932 11840 7984 11892
rect 8116 11883 8168 11892
rect 8116 11849 8125 11883
rect 8125 11849 8159 11883
rect 8159 11849 8168 11883
rect 8116 11840 8168 11849
rect 9128 11883 9180 11892
rect 9128 11849 9137 11883
rect 9137 11849 9171 11883
rect 9171 11849 9180 11883
rect 9128 11840 9180 11849
rect 7104 11772 7156 11824
rect 10692 11772 10744 11824
rect 15844 11772 15896 11824
rect 8944 11747 8996 11756
rect 8944 11713 8953 11747
rect 8953 11713 8987 11747
rect 8987 11713 8996 11747
rect 8944 11704 8996 11713
rect 9220 11747 9272 11756
rect 9220 11713 9229 11747
rect 9229 11713 9263 11747
rect 9263 11713 9272 11747
rect 9220 11704 9272 11713
rect 6276 11636 6328 11688
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 1860 11543 1912 11552
rect 1860 11509 1869 11543
rect 1869 11509 1903 11543
rect 1903 11509 1912 11543
rect 1860 11500 1912 11509
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 8300 11500 8352 11552
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 7566 11398 7618 11450
rect 7630 11398 7682 11450
rect 7694 11398 7746 11450
rect 7758 11398 7810 11450
rect 7822 11398 7874 11450
rect 3976 11296 4028 11348
rect 11152 11296 11204 11348
rect 11428 11296 11480 11348
rect 8208 11271 8260 11280
rect 8208 11237 8217 11271
rect 8217 11237 8251 11271
rect 8251 11237 8260 11271
rect 8208 11228 8260 11237
rect 9128 11271 9180 11280
rect 9128 11237 9137 11271
rect 9137 11237 9171 11271
rect 9171 11237 9180 11271
rect 9128 11228 9180 11237
rect 572 11160 624 11212
rect 4988 11203 5040 11212
rect 4988 11169 4997 11203
rect 4997 11169 5031 11203
rect 5031 11169 5040 11203
rect 4988 11160 5040 11169
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 1860 11092 1912 11144
rect 7196 11135 7248 11144
rect 2688 11024 2740 11076
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 5540 11067 5592 11076
rect 5540 11033 5549 11067
rect 5549 11033 5583 11067
rect 5583 11033 5592 11067
rect 5540 11024 5592 11033
rect 7288 11024 7340 11076
rect 8024 11024 8076 11076
rect 8484 11092 8536 11144
rect 16580 11092 16632 11144
rect 3148 10956 3200 11008
rect 9864 11024 9916 11076
rect 9220 10956 9272 11008
rect 16120 10956 16172 11008
rect 16580 10956 16632 11008
rect 3566 10854 3618 10906
rect 3630 10854 3682 10906
rect 3694 10854 3746 10906
rect 3758 10854 3810 10906
rect 3822 10854 3874 10906
rect 8566 10854 8618 10906
rect 8630 10854 8682 10906
rect 8694 10854 8746 10906
rect 8758 10854 8810 10906
rect 8822 10854 8874 10906
rect 15108 10888 15160 10940
rect 15476 10888 15528 10940
rect 16396 10888 16448 10940
rect 2228 10684 2280 10736
rect 4160 10684 4212 10736
rect 5632 10752 5684 10804
rect 7196 10684 7248 10736
rect 1768 10616 1820 10668
rect 2412 10616 2464 10668
rect 2780 10616 2832 10668
rect 5356 10616 5408 10668
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 6828 10616 6880 10668
rect 8208 10659 8260 10668
rect 8208 10625 8217 10659
rect 8217 10625 8251 10659
rect 8251 10625 8260 10659
rect 8208 10616 8260 10625
rect 1032 10548 1084 10600
rect 6368 10591 6420 10600
rect 6368 10557 6377 10591
rect 6377 10557 6411 10591
rect 6411 10557 6420 10591
rect 6368 10548 6420 10557
rect 8024 10480 8076 10532
rect 13452 10480 13504 10532
rect 14280 10480 14332 10532
rect 15568 10480 15620 10532
rect 2228 10412 2280 10464
rect 5356 10412 5408 10464
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9128 10412 9180 10421
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 7566 10310 7618 10362
rect 7630 10310 7682 10362
rect 7694 10310 7746 10362
rect 7758 10310 7810 10362
rect 7822 10310 7874 10362
rect 8944 10251 8996 10260
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 9220 10208 9272 10260
rect 15476 10208 15528 10260
rect 16396 10208 16448 10260
rect 3148 10072 3200 10124
rect 6000 10115 6052 10124
rect 6000 10081 6009 10115
rect 6009 10081 6043 10115
rect 6043 10081 6052 10115
rect 6000 10072 6052 10081
rect 9220 10072 9272 10124
rect 13912 10072 13964 10124
rect 14372 10072 14424 10124
rect 1492 10004 1544 10056
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 3056 10004 3108 10056
rect 5172 10004 5224 10056
rect 6460 10004 6512 10056
rect 9128 10004 9180 10056
rect 13728 10004 13780 10056
rect 16304 10004 16356 10056
rect 3240 9936 3292 9988
rect 7104 9936 7156 9988
rect 9312 9979 9364 9988
rect 9312 9945 9321 9979
rect 9321 9945 9355 9979
rect 9355 9945 9364 9979
rect 9312 9936 9364 9945
rect 16488 10072 16540 10124
rect 2320 9868 2372 9920
rect 3148 9868 3200 9920
rect 6644 9868 6696 9920
rect 6828 9868 6880 9920
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 8392 9868 8444 9920
rect 9404 9868 9456 9920
rect 3566 9766 3618 9818
rect 3630 9766 3682 9818
rect 3694 9766 3746 9818
rect 3758 9766 3810 9818
rect 3822 9766 3874 9818
rect 8566 9766 8618 9818
rect 8630 9766 8682 9818
rect 8694 9766 8746 9818
rect 8758 9766 8810 9818
rect 8822 9766 8874 9818
rect 1768 9664 1820 9716
rect 4896 9664 4948 9716
rect 1676 9596 1728 9648
rect 4620 9596 4672 9648
rect 2136 9528 2188 9580
rect 3424 9528 3476 9580
rect 5172 9528 5224 9580
rect 7012 9596 7064 9648
rect 9128 9639 9180 9648
rect 9128 9605 9137 9639
rect 9137 9605 9171 9639
rect 9171 9605 9180 9639
rect 9128 9596 9180 9605
rect 6828 9528 6880 9580
rect 4068 9460 4120 9512
rect 5816 9503 5868 9512
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 5816 9460 5868 9469
rect 13820 9460 13872 9512
rect 15384 9460 15436 9512
rect 848 9324 900 9376
rect 3884 9324 3936 9376
rect 6736 9367 6788 9376
rect 6736 9333 6745 9367
rect 6745 9333 6779 9367
rect 6779 9333 6788 9367
rect 6736 9324 6788 9333
rect 9036 9324 9088 9376
rect 15292 9324 15344 9376
rect 15568 9324 15620 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 7566 9222 7618 9274
rect 7630 9222 7682 9274
rect 7694 9222 7746 9274
rect 7758 9222 7810 9274
rect 7822 9222 7874 9274
rect 15568 9188 15620 9240
rect 15752 9188 15804 9240
rect 1584 9120 1636 9172
rect 2780 9120 2832 9172
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 4712 9163 4764 9172
rect 4712 9129 4721 9163
rect 4721 9129 4755 9163
rect 4755 9129 4764 9163
rect 4712 9120 4764 9129
rect 2872 9052 2924 9104
rect 3148 9052 3200 9104
rect 15752 9052 15804 9104
rect 16488 9800 16540 9852
rect 3056 8984 3108 9036
rect 3332 8984 3384 9036
rect 4160 8916 4212 8968
rect 5448 8916 5500 8968
rect 6552 8916 6604 8968
rect 9036 8959 9088 8968
rect 9036 8925 9045 8959
rect 9045 8925 9079 8959
rect 9079 8925 9088 8959
rect 9036 8916 9088 8925
rect 15384 8916 15436 8968
rect 15660 8916 15712 8968
rect 3424 8848 3476 8900
rect 7380 8848 7432 8900
rect 5540 8780 5592 8832
rect 6276 8780 6328 8832
rect 9128 8823 9180 8832
rect 9128 8789 9137 8823
rect 9137 8789 9171 8823
rect 9171 8789 9180 8823
rect 9128 8780 9180 8789
rect 15660 8780 15712 8832
rect 16488 8780 16540 8832
rect 3566 8678 3618 8730
rect 3630 8678 3682 8730
rect 3694 8678 3746 8730
rect 3758 8678 3810 8730
rect 3822 8678 3874 8730
rect 8566 8678 8618 8730
rect 8630 8678 8682 8730
rect 8694 8678 8746 8730
rect 8758 8678 8810 8730
rect 8822 8678 8874 8730
rect 16488 8644 16540 8696
rect 3240 8576 3292 8628
rect 6460 8576 6512 8628
rect 16580 8576 16632 8628
rect 4528 8508 4580 8560
rect 9128 8551 9180 8560
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 9128 8517 9137 8551
rect 9137 8517 9171 8551
rect 9171 8517 9180 8551
rect 9128 8508 9180 8517
rect 2872 8372 2924 8424
rect 5632 8440 5684 8492
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 15568 8440 15620 8492
rect 3792 8372 3844 8424
rect 6736 8372 6788 8424
rect 8208 8415 8260 8424
rect 8208 8381 8217 8415
rect 8217 8381 8251 8415
rect 8251 8381 8260 8415
rect 8208 8372 8260 8381
rect 9588 8372 9640 8424
rect 1768 8347 1820 8356
rect 1768 8313 1777 8347
rect 1777 8313 1811 8347
rect 1811 8313 1820 8347
rect 1768 8304 1820 8313
rect 2780 8304 2832 8356
rect 6828 8304 6880 8356
rect 1952 8236 2004 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 7566 8134 7618 8186
rect 7630 8134 7682 8186
rect 7694 8134 7746 8186
rect 7758 8134 7810 8186
rect 7822 8134 7874 8186
rect 2044 8032 2096 8084
rect 2964 8032 3016 8084
rect 4068 8032 4120 8084
rect 4252 7828 4304 7880
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 7012 7871 7064 7880
rect 4344 7828 4396 7837
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 8944 7871 8996 7880
rect 8944 7837 8953 7871
rect 8953 7837 8987 7871
rect 8987 7837 8996 7871
rect 8944 7828 8996 7837
rect 15476 7828 15528 7880
rect 16580 8440 16632 8492
rect 16672 8372 16724 8424
rect 16488 8236 16540 8288
rect 16580 8168 16632 8220
rect 9128 7803 9180 7812
rect 9128 7769 9137 7803
rect 9137 7769 9171 7803
rect 9171 7769 9180 7803
rect 9128 7760 9180 7769
rect 3700 7692 3752 7744
rect 4252 7692 4304 7744
rect 6276 7692 6328 7744
rect 7012 7692 7064 7744
rect 9404 7692 9456 7744
rect 3566 7590 3618 7642
rect 3630 7590 3682 7642
rect 3694 7590 3746 7642
rect 3758 7590 3810 7642
rect 3822 7590 3874 7642
rect 8566 7590 8618 7642
rect 8630 7590 8682 7642
rect 8694 7590 8746 7642
rect 8758 7590 8810 7642
rect 8822 7590 8874 7642
rect 5356 7488 5408 7540
rect 8024 7488 8076 7540
rect 8300 7488 8352 7540
rect 4068 7420 4120 7472
rect 4252 7420 4304 7472
rect 7104 7420 7156 7472
rect 1492 7352 1544 7404
rect 3056 7352 3108 7404
rect 8024 7352 8076 7404
rect 9772 7352 9824 7404
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 3056 7216 3108 7268
rect 3240 7216 3292 7268
rect 6368 7327 6420 7336
rect 6368 7293 6377 7327
rect 6377 7293 6411 7327
rect 6411 7293 6420 7327
rect 6368 7284 6420 7293
rect 6736 7327 6788 7336
rect 6736 7293 6745 7327
rect 6745 7293 6779 7327
rect 6779 7293 6788 7327
rect 6736 7284 6788 7293
rect 9772 7216 9824 7268
rect 16488 7216 16540 7268
rect 4160 7148 4212 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 7566 7046 7618 7098
rect 7630 7046 7682 7098
rect 7694 7046 7746 7098
rect 7758 7046 7810 7098
rect 7822 7046 7874 7098
rect 11336 7012 11388 7064
rect 16028 7012 16080 7064
rect 16580 7012 16632 7064
rect 1952 6944 2004 6996
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 3332 6808 3384 6860
rect 4344 6944 4396 6996
rect 4160 6876 4212 6928
rect 8300 6876 8352 6928
rect 8944 6876 8996 6928
rect 10600 6808 10652 6860
rect 15844 6808 15896 6860
rect 4252 6740 4304 6792
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 6092 6783 6144 6792
rect 5632 6740 5684 6749
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 8024 6740 8076 6792
rect 8300 6740 8352 6792
rect 7196 6672 7248 6724
rect 8944 6715 8996 6724
rect 8944 6681 8953 6715
rect 8953 6681 8987 6715
rect 8987 6681 8996 6715
rect 8944 6672 8996 6681
rect 9128 6715 9180 6724
rect 9128 6681 9137 6715
rect 9137 6681 9171 6715
rect 9171 6681 9180 6715
rect 9128 6672 9180 6681
rect 13268 6672 13320 6724
rect 16120 6672 16172 6724
rect 5540 6604 5592 6656
rect 9036 6604 9088 6656
rect 15844 6604 15896 6656
rect 16212 6604 16264 6656
rect 3566 6502 3618 6554
rect 3630 6502 3682 6554
rect 3694 6502 3746 6554
rect 3758 6502 3810 6554
rect 3822 6502 3874 6554
rect 8566 6502 8618 6554
rect 8630 6502 8682 6554
rect 8694 6502 8746 6554
rect 8758 6502 8810 6554
rect 8822 6502 8874 6554
rect 15476 6468 15528 6520
rect 16212 6468 16264 6520
rect 2228 6443 2280 6452
rect 2228 6409 2237 6443
rect 2237 6409 2271 6443
rect 2271 6409 2280 6443
rect 2228 6400 2280 6409
rect 3240 6400 3292 6452
rect 5816 6400 5868 6452
rect 4252 6332 4304 6384
rect 5356 6332 5408 6384
rect 7288 6400 7340 6452
rect 7472 6400 7524 6452
rect 9128 6400 9180 6452
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 2136 6264 2188 6316
rect 7380 6332 7432 6384
rect 7012 6307 7064 6316
rect 1492 6171 1544 6180
rect 1492 6137 1501 6171
rect 1501 6137 1535 6171
rect 1535 6137 1544 6171
rect 1492 6128 1544 6137
rect 4068 6060 4120 6112
rect 5632 6196 5684 6248
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 13820 6264 13872 6316
rect 6920 6196 6972 6248
rect 5632 6060 5684 6112
rect 8944 6103 8996 6112
rect 8944 6069 8953 6103
rect 8953 6069 8987 6103
rect 8987 6069 8996 6103
rect 8944 6060 8996 6069
rect 13912 6060 13964 6112
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 7566 5958 7618 6010
rect 7630 5958 7682 6010
rect 7694 5958 7746 6010
rect 7758 5958 7810 6010
rect 7822 5958 7874 6010
rect 13820 5992 13872 6044
rect 14372 5992 14424 6044
rect 16672 5992 16724 6044
rect 2964 5856 3016 5908
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 6184 5856 6236 5908
rect 9128 5899 9180 5908
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 3148 5788 3200 5840
rect 756 5720 808 5772
rect 2044 5652 2096 5704
rect 2228 5763 2280 5772
rect 2228 5729 2237 5763
rect 2237 5729 2271 5763
rect 2271 5729 2280 5763
rect 2228 5720 2280 5729
rect 4068 5720 4120 5772
rect 6828 5763 6880 5772
rect 6828 5729 6837 5763
rect 6837 5729 6871 5763
rect 6871 5729 6880 5763
rect 6828 5720 6880 5729
rect 8208 5763 8260 5772
rect 8208 5729 8217 5763
rect 8217 5729 8251 5763
rect 8251 5729 8260 5763
rect 8208 5720 8260 5729
rect 2780 5652 2832 5704
rect 3516 5652 3568 5704
rect 2688 5584 2740 5636
rect 3332 5584 3384 5636
rect 4344 5584 4396 5636
rect 8392 5652 8444 5704
rect 8208 5584 8260 5636
rect 5540 5516 5592 5568
rect 6828 5516 6880 5568
rect 7380 5516 7432 5568
rect 15752 5516 15804 5568
rect 3566 5414 3618 5466
rect 3630 5414 3682 5466
rect 3694 5414 3746 5466
rect 3758 5414 3810 5466
rect 3822 5414 3874 5466
rect 8566 5414 8618 5466
rect 8630 5414 8682 5466
rect 8694 5414 8746 5466
rect 8758 5414 8810 5466
rect 8822 5414 8874 5466
rect 13544 5448 13596 5500
rect 14188 5448 14240 5500
rect 4068 5312 4120 5364
rect 4896 5312 4948 5364
rect 6460 5312 6512 5364
rect 6736 5312 6788 5364
rect 572 5244 624 5296
rect 2780 5176 2832 5228
rect 5816 5244 5868 5296
rect 7288 5287 7340 5296
rect 7288 5253 7297 5287
rect 7297 5253 7331 5287
rect 7331 5253 7340 5287
rect 7288 5244 7340 5253
rect 7380 5244 7432 5296
rect 9312 5244 9364 5296
rect 4804 5176 4856 5228
rect 6184 5219 6236 5228
rect 6184 5185 6193 5219
rect 6193 5185 6227 5219
rect 6227 5185 6236 5219
rect 6184 5176 6236 5185
rect 6736 5176 6788 5228
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 8576 5176 8628 5228
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 4160 5108 4212 5160
rect 5540 5108 5592 5160
rect 7012 5108 7064 5160
rect 4528 5040 4580 5092
rect 4988 5040 5040 5092
rect 7472 4972 7524 5024
rect 8300 4972 8352 5024
rect 112 4836 164 4888
rect 2780 4836 2832 4888
rect 7566 4870 7618 4922
rect 7630 4870 7682 4922
rect 7694 4870 7746 4922
rect 7758 4870 7810 4922
rect 7822 4870 7874 4922
rect 1124 4768 1176 4820
rect 2412 4768 2464 4820
rect 5540 4768 5592 4820
rect 6092 4768 6144 4820
rect 6920 4768 6972 4820
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 940 4700 992 4752
rect 4160 4700 4212 4752
rect 1124 4632 1176 4684
rect 1308 4632 1360 4684
rect 3424 4632 3476 4684
rect 4896 4675 4948 4684
rect 1216 4564 1268 4616
rect 1860 4564 1912 4616
rect 2872 4564 2924 4616
rect 3700 4607 3752 4616
rect 3700 4573 3709 4607
rect 3709 4573 3743 4607
rect 3743 4573 3752 4607
rect 3700 4564 3752 4573
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 6644 4632 6696 4684
rect 8392 4632 8444 4684
rect 6276 4564 6328 4616
rect 8944 4564 8996 4616
rect 9312 4632 9364 4684
rect 4068 4496 4120 4548
rect 9312 4539 9364 4548
rect 9312 4505 9321 4539
rect 9321 4505 9355 4539
rect 9355 4505 9364 4539
rect 9312 4496 9364 4505
rect 4252 4428 4304 4480
rect 3566 4326 3618 4378
rect 3630 4326 3682 4378
rect 3694 4326 3746 4378
rect 3758 4326 3810 4378
rect 3822 4326 3874 4378
rect 8566 4326 8618 4378
rect 8630 4326 8682 4378
rect 8694 4326 8746 4378
rect 8758 4326 8810 4378
rect 8822 4326 8874 4378
rect 4436 4224 4488 4276
rect 8208 4224 8260 4276
rect 4160 4088 4212 4140
rect 4896 4088 4948 4140
rect 7012 4088 7064 4140
rect 8208 4088 8260 4140
rect 9220 4088 9272 4140
rect 12348 4088 12400 4140
rect 12440 4088 12492 4140
rect 4068 4063 4120 4072
rect 4068 4029 4077 4063
rect 4077 4029 4111 4063
rect 4111 4029 4120 4063
rect 4068 4020 4120 4029
rect 6552 4020 6604 4072
rect 6276 3995 6328 4004
rect 6276 3961 6285 3995
rect 6285 3961 6319 3995
rect 6319 3961 6328 3995
rect 6276 3952 6328 3961
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 7288 3884 7340 3936
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 7566 3782 7618 3834
rect 7630 3782 7682 3834
rect 7694 3782 7746 3834
rect 7758 3782 7810 3834
rect 7822 3782 7874 3834
rect 4620 3680 4672 3732
rect 5080 3680 5132 3732
rect 6092 3723 6144 3732
rect 6092 3689 6101 3723
rect 6101 3689 6135 3723
rect 6135 3689 6144 3723
rect 6092 3680 6144 3689
rect 6828 3723 6880 3732
rect 6828 3689 6837 3723
rect 6837 3689 6871 3723
rect 6871 3689 6880 3723
rect 6828 3680 6880 3689
rect 7196 3680 7248 3732
rect 8024 3723 8076 3732
rect 8024 3689 8033 3723
rect 8033 3689 8067 3723
rect 8067 3689 8076 3723
rect 8024 3680 8076 3689
rect 5172 3612 5224 3664
rect 6552 3544 6604 3596
rect 3516 3519 3568 3528
rect 3516 3485 3525 3519
rect 3525 3485 3559 3519
rect 3559 3485 3568 3519
rect 3516 3476 3568 3485
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4528 3476 4580 3528
rect 4712 3476 4764 3528
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 6644 3476 6696 3528
rect 8116 3476 8168 3528
rect 9404 3544 9456 3596
rect 9128 3476 9180 3528
rect 5080 3408 5132 3460
rect 5724 3408 5776 3460
rect 10324 3408 10376 3460
rect 16212 3408 16264 3460
rect 9220 3383 9272 3392
rect 9220 3349 9229 3383
rect 9229 3349 9263 3383
rect 9263 3349 9272 3383
rect 9220 3340 9272 3349
rect 3566 3238 3618 3290
rect 3630 3238 3682 3290
rect 3694 3238 3746 3290
rect 3758 3238 3810 3290
rect 3822 3238 3874 3290
rect 8566 3238 8618 3290
rect 8630 3238 8682 3290
rect 8694 3238 8746 3290
rect 8758 3238 8810 3290
rect 8822 3238 8874 3290
rect 3240 3136 3292 3188
rect 4988 3179 5040 3188
rect 4988 3145 4997 3179
rect 4997 3145 5031 3179
rect 5031 3145 5040 3179
rect 4988 3136 5040 3145
rect 6000 3136 6052 3188
rect 6736 3136 6788 3188
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 8484 3136 8536 3188
rect 9220 3179 9272 3188
rect 9220 3145 9229 3179
rect 9229 3145 9263 3179
rect 9263 3145 9272 3179
rect 9220 3136 9272 3145
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 4252 3000 4304 3052
rect 5632 3068 5684 3120
rect 4436 3000 4488 3052
rect 4896 3043 4948 3052
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 13912 3068 13964 3120
rect 7472 3000 7524 3052
rect 9772 3000 9824 3052
rect 14096 2864 14148 2916
rect 16396 2864 16448 2916
rect 3884 2796 3936 2848
rect 7566 2694 7618 2746
rect 7630 2694 7682 2746
rect 7694 2694 7746 2746
rect 7758 2694 7810 2746
rect 7822 2694 7874 2746
rect 4160 2592 4212 2644
rect 8024 2592 8076 2644
rect 9036 2592 9088 2644
rect 2780 2456 2832 2508
rect 4528 2388 4580 2440
rect 5080 2388 5132 2440
rect 7380 2456 7432 2508
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 9404 2456 9456 2508
rect 8484 2388 8536 2440
rect 9956 2388 10008 2440
rect 3148 2252 3200 2304
rect 4896 2295 4948 2304
rect 4896 2261 4905 2295
rect 4905 2261 4939 2295
rect 4939 2261 4948 2295
rect 4896 2252 4948 2261
rect 6000 2295 6052 2304
rect 6000 2261 6009 2295
rect 6009 2261 6043 2295
rect 6043 2261 6052 2295
rect 6000 2252 6052 2261
rect 8116 2252 8168 2304
rect 3566 2150 3618 2202
rect 3630 2150 3682 2202
rect 3694 2150 3746 2202
rect 3758 2150 3810 2202
rect 3822 2150 3874 2202
rect 8566 2150 8618 2202
rect 8630 2150 8682 2202
rect 8694 2150 8746 2202
rect 8758 2150 8810 2202
rect 8822 2150 8874 2202
rect 3332 2048 3384 2100
rect 4068 1980 4120 2032
rect 3976 1912 4028 1964
rect 5448 2048 5500 2100
rect 5632 2091 5684 2100
rect 5632 2057 5641 2091
rect 5641 2057 5675 2091
rect 5675 2057 5684 2091
rect 5632 2048 5684 2057
rect 8484 2048 8536 2100
rect 9496 2048 9548 2100
rect 4344 1980 4396 2032
rect 6000 1980 6052 2032
rect 4804 1955 4856 1964
rect 4804 1921 4813 1955
rect 4813 1921 4847 1955
rect 4847 1921 4856 1955
rect 4804 1912 4856 1921
rect 5080 1912 5132 1964
rect 5448 1955 5500 1964
rect 5448 1921 5457 1955
rect 5457 1921 5491 1955
rect 5491 1921 5500 1955
rect 5448 1912 5500 1921
rect 6092 1955 6144 1964
rect 6092 1921 6101 1955
rect 6101 1921 6135 1955
rect 6135 1921 6144 1955
rect 6092 1912 6144 1921
rect 9036 1980 9088 2032
rect 6920 1955 6972 1964
rect 6920 1921 6929 1955
rect 6929 1921 6963 1955
rect 6963 1921 6972 1955
rect 6920 1912 6972 1921
rect 9220 1912 9272 1964
rect 9588 1912 9640 1964
rect 4252 1819 4304 1828
rect 4252 1785 4261 1819
rect 4261 1785 4295 1819
rect 4295 1785 4304 1819
rect 4252 1776 4304 1785
rect 6276 1751 6328 1760
rect 6276 1717 6285 1751
rect 6285 1717 6319 1751
rect 6319 1717 6328 1751
rect 6276 1708 6328 1717
rect 6828 1751 6880 1760
rect 6828 1717 6837 1751
rect 6837 1717 6871 1751
rect 6871 1717 6880 1751
rect 6828 1708 6880 1717
rect 7566 1606 7618 1658
rect 7630 1606 7682 1658
rect 7694 1606 7746 1658
rect 7758 1606 7810 1658
rect 7822 1606 7874 1658
rect 16672 5516 16724 5568
rect 16672 1572 16724 1624
rect 664 1504 716 1556
rect 4896 1504 4948 1556
rect 204 1436 256 1488
rect 4804 1436 4856 1488
rect 8944 1479 8996 1488
rect 8944 1445 8953 1479
rect 8953 1445 8987 1479
rect 8987 1445 8996 1479
rect 8944 1436 8996 1445
rect 388 1368 440 1420
rect 5448 1368 5500 1420
rect 6828 1368 6880 1420
rect 2964 1300 3016 1352
rect 4436 1300 4488 1352
rect 4804 1343 4856 1352
rect 4804 1309 4813 1343
rect 4813 1309 4847 1343
rect 4847 1309 4856 1343
rect 4804 1300 4856 1309
rect 5080 1300 5132 1352
rect 5264 1300 5316 1352
rect 6736 1343 6788 1352
rect 4252 1275 4304 1284
rect 4252 1241 4261 1275
rect 4261 1241 4295 1275
rect 4295 1241 4304 1275
rect 4252 1232 4304 1241
rect 6736 1309 6745 1343
rect 6745 1309 6779 1343
rect 6779 1309 6788 1343
rect 6736 1300 6788 1309
rect 8208 1300 8260 1352
rect 4068 1164 4120 1216
rect 4988 1207 5040 1216
rect 4988 1173 4997 1207
rect 4997 1173 5031 1207
rect 5031 1173 5040 1207
rect 4988 1164 5040 1173
rect 6092 1207 6144 1216
rect 6092 1173 6101 1207
rect 6101 1173 6135 1207
rect 6135 1173 6144 1207
rect 6092 1164 6144 1173
rect 6552 1207 6604 1216
rect 6552 1173 6561 1207
rect 6561 1173 6595 1207
rect 6595 1173 6604 1207
rect 6552 1164 6604 1173
rect 7380 1207 7432 1216
rect 7380 1173 7389 1207
rect 7389 1173 7423 1207
rect 7423 1173 7432 1207
rect 7380 1164 7432 1173
rect 9128 1207 9180 1216
rect 9128 1173 9137 1207
rect 9137 1173 9171 1207
rect 9171 1173 9180 1207
rect 9128 1164 9180 1173
rect 3566 1062 3618 1114
rect 3630 1062 3682 1114
rect 3694 1062 3746 1114
rect 3758 1062 3810 1114
rect 3822 1062 3874 1114
rect 8566 1062 8618 1114
rect 8630 1062 8682 1114
rect 8694 1062 8746 1114
rect 8758 1062 8810 1114
rect 8822 1062 8874 1114
<< metal2 >>
rect 492 16238 888 16266
rect 386 15464 442 15473
rect 386 15399 442 15408
rect 296 14884 348 14890
rect 296 14826 348 14832
rect 112 12640 164 12646
rect 112 12582 164 12588
rect 124 4894 152 12582
rect 202 10704 258 10713
rect 202 10639 258 10648
rect 112 4888 164 4894
rect 112 4830 164 4836
rect 216 1494 244 10639
rect 204 1488 256 1494
rect 204 1430 256 1436
rect 308 785 336 14826
rect 400 1426 428 15399
rect 492 15094 520 16238
rect 860 16130 888 16238
rect 938 16200 994 17000
rect 1398 16200 1454 17000
rect 1858 16200 1914 17000
rect 2318 16200 2374 17000
rect 2778 16200 2834 17000
rect 2884 16238 3096 16266
rect 952 16130 980 16200
rect 860 16102 980 16130
rect 1412 15434 1440 16200
rect 1400 15428 1452 15434
rect 1400 15370 1452 15376
rect 1216 15360 1268 15366
rect 1216 15302 1268 15308
rect 480 15088 532 15094
rect 480 15030 532 15036
rect 492 1601 520 15030
rect 756 14612 808 14618
rect 756 14554 808 14560
rect 662 13968 718 13977
rect 662 13903 718 13912
rect 572 11212 624 11218
rect 572 11154 624 11160
rect 584 5302 612 11154
rect 572 5296 624 5302
rect 572 5238 624 5244
rect 478 1592 534 1601
rect 676 1562 704 13903
rect 768 5778 796 14554
rect 1122 13288 1178 13297
rect 1122 13223 1178 13232
rect 940 13184 992 13190
rect 940 13126 992 13132
rect 848 9376 900 9382
rect 848 9318 900 9324
rect 756 5772 808 5778
rect 756 5714 808 5720
rect 478 1527 534 1536
rect 664 1556 716 1562
rect 664 1498 716 1504
rect 388 1420 440 1426
rect 388 1362 440 1368
rect 860 1193 888 9318
rect 952 4758 980 13126
rect 1032 10600 1084 10606
rect 1032 10542 1084 10548
rect 940 4752 992 4758
rect 940 4694 992 4700
rect 1044 1465 1072 10542
rect 1136 4826 1164 13223
rect 1124 4820 1176 4826
rect 1124 4762 1176 4768
rect 1124 4684 1176 4690
rect 1124 4626 1176 4632
rect 1030 1456 1086 1465
rect 1030 1391 1086 1400
rect 1136 1329 1164 4626
rect 1228 4622 1256 15302
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1308 13932 1360 13938
rect 1308 13874 1360 13880
rect 1320 4690 1348 13874
rect 1504 12889 1532 14758
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1596 13870 1624 14214
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1582 13016 1638 13025
rect 1582 12951 1638 12960
rect 1490 12880 1546 12889
rect 1596 12850 1624 12951
rect 1490 12815 1546 12824
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1596 12186 1624 12786
rect 1872 12458 1900 16200
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1504 12158 1624 12186
rect 1688 12430 1900 12458
rect 1504 10062 1532 12158
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1596 11150 1624 12038
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1596 9178 1624 11086
rect 1688 9654 1716 12430
rect 2056 12102 2084 13806
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11150 1900 11494
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1780 10062 1808 10610
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1780 9722 1808 9998
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1950 9616 2006 9625
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 6866 1532 7346
rect 1688 6914 1716 9590
rect 2148 9586 2176 15370
rect 2332 13410 2360 16200
rect 2792 16130 2820 16200
rect 2884 16130 2912 16238
rect 2792 16102 2912 16130
rect 2566 15804 2874 15813
rect 2566 15802 2572 15804
rect 2628 15802 2652 15804
rect 2708 15802 2732 15804
rect 2788 15802 2812 15804
rect 2868 15802 2874 15804
rect 2628 15750 2630 15802
rect 2810 15750 2812 15802
rect 2566 15748 2572 15750
rect 2628 15748 2652 15750
rect 2708 15748 2732 15750
rect 2788 15748 2812 15750
rect 2868 15748 2874 15750
rect 2566 15739 2874 15748
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2700 15178 2728 15438
rect 2700 15150 2820 15178
rect 2792 14890 2820 15150
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2566 14716 2874 14725
rect 2566 14714 2572 14716
rect 2628 14714 2652 14716
rect 2708 14714 2732 14716
rect 2788 14714 2812 14716
rect 2868 14714 2874 14716
rect 2628 14662 2630 14714
rect 2810 14662 2812 14714
rect 2566 14660 2572 14662
rect 2628 14660 2652 14662
rect 2708 14660 2732 14662
rect 2788 14660 2812 14662
rect 2868 14660 2874 14662
rect 2566 14651 2874 14660
rect 2504 14340 2556 14346
rect 2504 14282 2556 14288
rect 2412 13864 2464 13870
rect 2516 13841 2544 14282
rect 2412 13806 2464 13812
rect 2502 13832 2558 13841
rect 2240 13382 2360 13410
rect 2240 10742 2268 13382
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2332 12209 2360 13194
rect 2424 12850 2452 13806
rect 2502 13767 2558 13776
rect 2566 13628 2874 13637
rect 2566 13626 2572 13628
rect 2628 13626 2652 13628
rect 2708 13626 2732 13628
rect 2788 13626 2812 13628
rect 2868 13626 2874 13628
rect 2628 13574 2630 13626
rect 2810 13574 2812 13626
rect 2566 13572 2572 13574
rect 2628 13572 2652 13574
rect 2708 13572 2732 13574
rect 2788 13572 2812 13574
rect 2868 13572 2874 13574
rect 2566 13563 2874 13572
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2504 12776 2556 12782
rect 2502 12744 2504 12753
rect 2556 12744 2558 12753
rect 2502 12679 2558 12688
rect 2566 12540 2874 12549
rect 2566 12538 2572 12540
rect 2628 12538 2652 12540
rect 2708 12538 2732 12540
rect 2788 12538 2812 12540
rect 2868 12538 2874 12540
rect 2628 12486 2630 12538
rect 2810 12486 2812 12538
rect 2566 12484 2572 12486
rect 2628 12484 2652 12486
rect 2708 12484 2732 12486
rect 2788 12484 2812 12486
rect 2868 12484 2874 12486
rect 2566 12475 2874 12484
rect 2686 12336 2742 12345
rect 2976 12306 3004 14894
rect 3068 13025 3096 16238
rect 3238 16200 3294 17000
rect 3698 16200 3754 17000
rect 4066 16552 4122 16561
rect 4066 16487 4122 16496
rect 3804 16238 4016 16266
rect 3252 15910 3280 16200
rect 3712 16130 3740 16200
rect 3804 16130 3832 16238
rect 3712 16102 3832 16130
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 3160 15026 3188 15370
rect 3566 15260 3874 15269
rect 3566 15258 3572 15260
rect 3628 15258 3652 15260
rect 3708 15258 3732 15260
rect 3788 15258 3812 15260
rect 3868 15258 3874 15260
rect 3628 15206 3630 15258
rect 3810 15206 3812 15258
rect 3566 15204 3572 15206
rect 3628 15204 3652 15206
rect 3708 15204 3732 15206
rect 3788 15204 3812 15206
rect 3868 15204 3874 15206
rect 3566 15195 3874 15204
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3160 14278 3188 14962
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3252 14482 3280 14826
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 3252 13852 3280 14418
rect 3896 14385 3924 14758
rect 3882 14376 3938 14385
rect 3882 14311 3938 14320
rect 3566 14172 3874 14181
rect 3566 14170 3572 14172
rect 3628 14170 3652 14172
rect 3708 14170 3732 14172
rect 3788 14170 3812 14172
rect 3868 14170 3874 14172
rect 3628 14118 3630 14170
rect 3810 14118 3812 14170
rect 3566 14116 3572 14118
rect 3628 14116 3652 14118
rect 3708 14116 3732 14118
rect 3788 14116 3812 14118
rect 3868 14116 3874 14118
rect 3566 14107 3874 14116
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3332 14000 3384 14006
rect 3330 13968 3332 13977
rect 3384 13968 3386 13977
rect 3330 13903 3386 13912
rect 3620 13870 3648 14010
rect 3608 13864 3660 13870
rect 3252 13824 3372 13852
rect 3238 13696 3294 13705
rect 3238 13631 3294 13640
rect 3252 13326 3280 13631
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3054 13016 3110 13025
rect 3054 12951 3110 12960
rect 3252 12481 3280 13262
rect 3238 12472 3294 12481
rect 3238 12407 3294 12416
rect 2686 12271 2742 12280
rect 2964 12300 3016 12306
rect 2318 12200 2374 12209
rect 2700 12170 2728 12271
rect 2964 12242 3016 12248
rect 2318 12135 2374 12144
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2700 11830 2728 12106
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2566 11452 2874 11461
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11387 2874 11396
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2228 10736 2280 10742
rect 2226 10704 2228 10713
rect 2280 10704 2282 10713
rect 2226 10639 2282 10648
rect 2410 10704 2466 10713
rect 2700 10690 2728 11018
rect 2700 10674 2820 10690
rect 2700 10668 2832 10674
rect 2700 10662 2780 10668
rect 2410 10639 2412 10648
rect 2464 10639 2466 10648
rect 2412 10610 2464 10616
rect 2780 10610 2832 10616
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 1950 9551 2006 9560
rect 2136 9580 2188 9586
rect 1964 8498 1992 9551
rect 2136 9522 2188 9528
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1766 8392 1822 8401
rect 1766 8327 1768 8336
rect 1820 8327 1822 8336
rect 1768 8298 1820 8304
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1964 7002 1992 8230
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1688 6886 1900 6914
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1490 6216 1546 6225
rect 1490 6151 1492 6160
rect 1544 6151 1546 6160
rect 1492 6122 1544 6128
rect 1688 4729 1716 6258
rect 1674 4720 1730 4729
rect 1308 4684 1360 4690
rect 1674 4655 1730 4664
rect 1308 4626 1360 4632
rect 1872 4622 1900 6886
rect 2056 5710 2084 8026
rect 2134 7848 2190 7857
rect 2134 7783 2190 7792
rect 2148 6322 2176 7783
rect 2240 6914 2268 10406
rect 2566 10364 2874 10373
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10299 2874 10308
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2332 7018 2360 9862
rect 2566 9276 2874 9285
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9211 2874 9220
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2792 8362 2820 9114
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2884 8430 2912 9046
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2566 8188 2874 8197
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8123 2874 8132
rect 2976 8090 3004 12242
rect 3344 12238 3372 13824
rect 3608 13806 3660 13812
rect 3566 13084 3874 13093
rect 3566 13082 3572 13084
rect 3628 13082 3652 13084
rect 3708 13082 3732 13084
rect 3788 13082 3812 13084
rect 3868 13082 3874 13084
rect 3628 13030 3630 13082
rect 3810 13030 3812 13082
rect 3566 13028 3572 13030
rect 3628 13028 3652 13030
rect 3708 13028 3732 13030
rect 3788 13028 3812 13030
rect 3868 13028 3874 13030
rect 3566 13019 3874 13028
rect 3884 12912 3936 12918
rect 3422 12880 3478 12889
rect 3422 12815 3478 12824
rect 3882 12880 3884 12889
rect 3936 12880 3938 12889
rect 3882 12815 3938 12824
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3344 11830 3372 12174
rect 3332 11824 3384 11830
rect 3332 11766 3384 11772
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10130 3188 10950
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3068 9042 3096 9998
rect 3240 9988 3292 9994
rect 3240 9930 3292 9936
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3160 9110 3188 9862
rect 3252 9178 3280 9930
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3344 9042 3372 11630
rect 3436 9586 3464 12815
rect 3988 12594 4016 16238
rect 4080 15706 4108 16487
rect 4158 16200 4214 17000
rect 4264 16238 4568 16266
rect 4172 16130 4200 16200
rect 4264 16130 4292 16238
rect 4172 16102 4292 16130
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4080 15201 4108 15438
rect 4158 15328 4214 15337
rect 4158 15263 4214 15272
rect 4066 15192 4122 15201
rect 4066 15127 4122 15136
rect 4080 15094 4108 15127
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 4172 14498 4200 15263
rect 4434 15056 4490 15065
rect 4434 14991 4490 15000
rect 4252 14952 4304 14958
rect 4344 14952 4396 14958
rect 4252 14894 4304 14900
rect 4342 14920 4344 14929
rect 4396 14920 4398 14929
rect 4080 14482 4200 14498
rect 4068 14476 4200 14482
rect 4120 14470 4200 14476
rect 4068 14418 4120 14424
rect 4068 14272 4120 14278
rect 4264 14249 4292 14894
rect 4342 14855 4398 14864
rect 4250 14240 4306 14249
rect 4120 14220 4200 14226
rect 4068 14214 4200 14220
rect 4080 14198 4200 14214
rect 4172 13394 4200 14198
rect 4250 14175 4306 14184
rect 4448 13938 4476 14991
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4540 13433 4568 16238
rect 4618 16200 4674 17000
rect 5078 16200 5134 17000
rect 5538 16200 5594 17000
rect 5998 16200 6054 17000
rect 6458 16200 6514 17000
rect 14186 16552 14242 16561
rect 14186 16487 14242 16496
rect 16670 16552 16726 16561
rect 16670 16487 16726 16496
rect 4632 15586 4660 16200
rect 4632 15558 4752 15586
rect 4618 15464 4674 15473
rect 4618 15399 4620 15408
rect 4672 15399 4674 15408
rect 4620 15370 4672 15376
rect 4724 13802 4752 15558
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4816 14074 4844 14826
rect 5092 14249 5120 16200
rect 5446 16144 5502 16153
rect 5446 16079 5502 16088
rect 5460 15570 5488 16079
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5552 15450 5580 16200
rect 5724 15496 5776 15502
rect 5552 15422 5672 15450
rect 5724 15438 5776 15444
rect 5540 15360 5592 15366
rect 5368 15308 5540 15314
rect 5368 15302 5592 15308
rect 5368 15286 5580 15302
rect 5368 14958 5396 15286
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5368 14346 5396 14894
rect 5644 14498 5672 15422
rect 5736 15162 5764 15438
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5460 14482 5672 14498
rect 5448 14476 5672 14482
rect 5500 14470 5672 14476
rect 5448 14418 5500 14424
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5540 14272 5592 14278
rect 5078 14240 5134 14249
rect 5540 14214 5592 14220
rect 5078 14175 5134 14184
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 4896 13864 4948 13870
rect 4894 13832 4896 13841
rect 4948 13832 4950 13841
rect 4712 13796 4764 13802
rect 4894 13767 4950 13776
rect 4712 13738 4764 13744
rect 4526 13424 4582 13433
rect 4160 13388 4212 13394
rect 4526 13359 4582 13368
rect 4160 13330 4212 13336
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 3988 12566 4200 12594
rect 4066 12472 4122 12481
rect 4066 12407 4122 12416
rect 4080 12345 4108 12407
rect 4066 12336 4122 12345
rect 4066 12271 4122 12280
rect 4068 12096 4120 12102
rect 3974 12064 4030 12073
rect 4068 12038 4120 12044
rect 3566 11996 3874 12005
rect 3974 11999 4030 12008
rect 3566 11994 3572 11996
rect 3628 11994 3652 11996
rect 3708 11994 3732 11996
rect 3788 11994 3812 11996
rect 3868 11994 3874 11996
rect 3628 11942 3630 11994
rect 3810 11942 3812 11994
rect 3566 11940 3572 11942
rect 3628 11940 3652 11942
rect 3708 11940 3732 11942
rect 3788 11940 3812 11942
rect 3868 11940 3874 11942
rect 3566 11931 3874 11940
rect 3988 11354 4016 11999
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3566 10908 3874 10917
rect 3566 10906 3572 10908
rect 3628 10906 3652 10908
rect 3708 10906 3732 10908
rect 3788 10906 3812 10908
rect 3868 10906 3874 10908
rect 3628 10854 3630 10906
rect 3810 10854 3812 10906
rect 3566 10852 3572 10854
rect 3628 10852 3652 10854
rect 3708 10852 3732 10854
rect 3788 10852 3812 10854
rect 3868 10852 3874 10854
rect 3566 10843 3874 10852
rect 4080 10169 4108 12038
rect 4172 11257 4200 12566
rect 4356 12481 4384 12786
rect 4342 12472 4398 12481
rect 4342 12407 4398 12416
rect 4724 12322 4752 13738
rect 5276 13394 5304 13942
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5172 13320 5224 13326
rect 5170 13288 5172 13297
rect 5224 13288 5226 13297
rect 5170 13223 5226 13232
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4816 12434 4844 12582
rect 4816 12406 4936 12434
rect 4724 12294 4844 12322
rect 4436 12232 4488 12238
rect 4342 12200 4398 12209
rect 4436 12174 4488 12180
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4342 12135 4398 12144
rect 4356 11558 4384 12135
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4158 11248 4214 11257
rect 4158 11183 4214 11192
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4066 10160 4122 10169
rect 4066 10095 4122 10104
rect 3566 9820 3874 9829
rect 3566 9818 3572 9820
rect 3628 9818 3652 9820
rect 3708 9818 3732 9820
rect 3788 9818 3812 9820
rect 3868 9818 3874 9820
rect 3628 9766 3630 9818
rect 3810 9766 3812 9818
rect 3566 9764 3572 9766
rect 3628 9764 3652 9766
rect 3708 9764 3732 9766
rect 3788 9764 3812 9766
rect 3868 9764 3874 9766
rect 3566 9755 3874 9764
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 3068 7410 3096 8978
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3146 8528 3202 8537
rect 3146 8463 3202 8472
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 2566 7100 2874 7109
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7035 2874 7044
rect 2962 7032 3018 7041
rect 2332 6990 2452 7018
rect 2240 6886 2360 6914
rect 2226 6488 2282 6497
rect 2226 6423 2228 6432
rect 2280 6423 2282 6432
rect 2228 6394 2280 6400
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2226 5808 2282 5817
rect 2226 5743 2228 5752
rect 2280 5743 2282 5752
rect 2228 5714 2280 5720
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 1216 4616 1268 4622
rect 1216 4558 1268 4564
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 2332 3074 2360 6886
rect 2424 5250 2452 6990
rect 2962 6967 3018 6976
rect 2566 6012 2874 6021
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5947 2874 5956
rect 2976 5914 3004 6967
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2780 5704 2832 5710
rect 2594 5672 2650 5681
rect 2780 5646 2832 5652
rect 2594 5607 2650 5616
rect 2688 5636 2740 5642
rect 2424 5222 2544 5250
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2424 3913 2452 4762
rect 2516 4049 2544 5222
rect 2502 4040 2558 4049
rect 2502 3975 2558 3984
rect 2410 3904 2466 3913
rect 2410 3839 2466 3848
rect 2608 3777 2636 5607
rect 2688 5578 2740 5584
rect 2594 3768 2650 3777
rect 2594 3703 2650 3712
rect 2410 3088 2466 3097
rect 2332 3046 2410 3074
rect 2410 3023 2466 3032
rect 2700 2496 2728 5578
rect 2792 5234 2820 5646
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2780 4888 2832 4894
rect 2780 4830 2832 4836
rect 2792 3777 2820 4830
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2778 3768 2834 3777
rect 2778 3703 2834 3712
rect 2884 3505 2912 4558
rect 3068 4185 3096 7210
rect 3160 5846 3188 8463
rect 3252 7274 3280 8570
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3344 7018 3372 8978
rect 3896 8922 3924 9318
rect 3424 8900 3476 8906
rect 3896 8894 4016 8922
rect 3424 8842 3476 8848
rect 3436 8514 3464 8842
rect 3566 8732 3874 8741
rect 3566 8730 3572 8732
rect 3628 8730 3652 8732
rect 3708 8730 3732 8732
rect 3788 8730 3812 8732
rect 3868 8730 3874 8732
rect 3628 8678 3630 8730
rect 3810 8678 3812 8730
rect 3566 8676 3572 8678
rect 3628 8676 3652 8678
rect 3708 8676 3732 8678
rect 3788 8676 3812 8678
rect 3868 8676 3874 8678
rect 3566 8667 3874 8676
rect 3988 8673 4016 8894
rect 3974 8664 4030 8673
rect 3974 8599 4030 8608
rect 3436 8486 3740 8514
rect 3422 8392 3478 8401
rect 3422 8327 3478 8336
rect 3252 6990 3372 7018
rect 3252 6458 3280 6990
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3238 5944 3294 5953
rect 3238 5879 3294 5888
rect 3148 5840 3200 5846
rect 3148 5782 3200 5788
rect 3146 4584 3202 4593
rect 3146 4519 3202 4528
rect 3054 4176 3110 4185
rect 3054 4111 3110 4120
rect 2870 3496 2926 3505
rect 2870 3431 2926 3440
rect 3160 2774 3188 4519
rect 3252 3194 3280 5879
rect 3344 5642 3372 6802
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3330 4720 3386 4729
rect 3436 4690 3464 8327
rect 3712 7750 3740 8486
rect 3792 8424 3844 8430
rect 3844 8372 4016 8378
rect 3792 8366 4016 8372
rect 3804 8350 4016 8366
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3566 7644 3874 7653
rect 3566 7642 3572 7644
rect 3628 7642 3652 7644
rect 3708 7642 3732 7644
rect 3788 7642 3812 7644
rect 3868 7642 3874 7644
rect 3628 7590 3630 7642
rect 3810 7590 3812 7642
rect 3566 7588 3572 7590
rect 3628 7588 3652 7590
rect 3708 7588 3732 7590
rect 3788 7588 3812 7590
rect 3868 7588 3874 7590
rect 3566 7579 3874 7588
rect 3566 6556 3874 6565
rect 3566 6554 3572 6556
rect 3628 6554 3652 6556
rect 3708 6554 3732 6556
rect 3788 6554 3812 6556
rect 3868 6554 3874 6556
rect 3628 6502 3630 6554
rect 3810 6502 3812 6554
rect 3566 6500 3572 6502
rect 3628 6500 3652 6502
rect 3708 6500 3732 6502
rect 3788 6500 3812 6502
rect 3868 6500 3874 6502
rect 3566 6491 3874 6500
rect 3516 5704 3568 5710
rect 3514 5672 3516 5681
rect 3568 5672 3570 5681
rect 3514 5607 3570 5616
rect 3566 5468 3874 5477
rect 3566 5466 3572 5468
rect 3628 5466 3652 5468
rect 3708 5466 3732 5468
rect 3788 5466 3812 5468
rect 3868 5466 3874 5468
rect 3628 5414 3630 5466
rect 3810 5414 3812 5466
rect 3566 5412 3572 5414
rect 3628 5412 3652 5414
rect 3708 5412 3732 5414
rect 3788 5412 3812 5414
rect 3868 5412 3874 5414
rect 3566 5403 3874 5412
rect 3698 5128 3754 5137
rect 3698 5063 3754 5072
rect 3330 4655 3386 4664
rect 3424 4684 3476 4690
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3344 2961 3372 4655
rect 3424 4626 3476 4632
rect 3712 4622 3740 5063
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3566 4380 3874 4389
rect 3566 4378 3572 4380
rect 3628 4378 3652 4380
rect 3708 4378 3732 4380
rect 3788 4378 3812 4380
rect 3868 4378 3874 4380
rect 3628 4326 3630 4378
rect 3810 4326 3812 4378
rect 3566 4324 3572 4326
rect 3628 4324 3652 4326
rect 3708 4324 3732 4326
rect 3788 4324 3812 4326
rect 3868 4324 3874 4326
rect 3566 4315 3874 4324
rect 3514 4040 3570 4049
rect 3514 3975 3570 3984
rect 3528 3534 3556 3975
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3566 3292 3874 3301
rect 3566 3290 3572 3292
rect 3628 3290 3652 3292
rect 3708 3290 3732 3292
rect 3788 3290 3812 3292
rect 3868 3290 3874 3292
rect 3628 3238 3630 3290
rect 3810 3238 3812 3290
rect 3566 3236 3572 3238
rect 3628 3236 3652 3238
rect 3708 3236 3732 3238
rect 3788 3236 3812 3238
rect 3868 3236 3874 3238
rect 3566 3227 3874 3236
rect 3514 3088 3570 3097
rect 3514 3023 3516 3032
rect 3568 3023 3570 3032
rect 3516 2994 3568 3000
rect 3330 2952 3386 2961
rect 3330 2887 3386 2896
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3160 2746 3372 2774
rect 2780 2508 2832 2514
rect 2700 2468 2780 2496
rect 2780 2450 2832 2456
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 1858 1592 1914 1601
rect 2318 1592 2374 1601
rect 1914 1550 2318 1578
rect 1858 1527 1914 1536
rect 2318 1527 2374 1536
rect 3160 1465 3188 2246
rect 3344 2106 3372 2746
rect 3896 2394 3924 2790
rect 3988 2774 4016 8350
rect 4080 8090 4108 9454
rect 4172 9081 4200 10678
rect 4356 9466 4384 11494
rect 4264 9438 4384 9466
rect 4158 9072 4214 9081
rect 4158 9007 4214 9016
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4172 7562 4200 8910
rect 4264 7886 4292 9438
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4080 7534 4200 7562
rect 4080 7478 4108 7534
rect 4264 7478 4292 7686
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 4080 6118 4108 7278
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4172 6934 4200 7142
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5778 4108 6054
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4066 5536 4122 5545
rect 4066 5471 4122 5480
rect 4080 5370 4108 5471
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4172 5166 4200 6870
rect 4264 6798 4292 7414
rect 4356 7002 4384 7822
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4264 6390 4292 6734
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 4264 5624 4292 6326
rect 4344 5636 4396 5642
rect 4264 5596 4344 5624
rect 4344 5578 4396 5584
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4066 4992 4122 5001
rect 4066 4927 4122 4936
rect 4080 4554 4108 4927
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 4172 4146 4200 4694
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4068 4072 4120 4078
rect 4066 4040 4068 4049
rect 4120 4040 4122 4049
rect 4066 3975 4122 3984
rect 4158 3768 4214 3777
rect 4158 3703 4214 3712
rect 4172 3534 4200 3703
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4264 3058 4292 4422
rect 4448 4282 4476 12174
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 4540 5953 4568 8502
rect 4526 5944 4582 5953
rect 4526 5879 4582 5888
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4342 4176 4398 4185
rect 4342 4111 4398 4120
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 3988 2746 4200 2774
rect 4066 2680 4122 2689
rect 4172 2650 4200 2746
rect 4066 2615 4122 2624
rect 4160 2644 4212 2650
rect 3896 2366 4016 2394
rect 3566 2204 3874 2213
rect 3566 2202 3572 2204
rect 3628 2202 3652 2204
rect 3708 2202 3732 2204
rect 3788 2202 3812 2204
rect 3868 2202 3874 2204
rect 3628 2150 3630 2202
rect 3810 2150 3812 2202
rect 3566 2148 3572 2150
rect 3628 2148 3652 2150
rect 3708 2148 3732 2150
rect 3788 2148 3812 2150
rect 3868 2148 3874 2150
rect 3566 2139 3874 2148
rect 3332 2100 3384 2106
rect 3332 2042 3384 2048
rect 3988 1970 4016 2366
rect 4080 2038 4108 2615
rect 4160 2586 4212 2592
rect 4356 2038 4384 4111
rect 4540 3534 4568 5034
rect 4632 3738 4660 9590
rect 4724 9178 4752 12174
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4816 9058 4844 12294
rect 4908 9722 4936 12406
rect 4986 12200 5042 12209
rect 4986 12135 5042 12144
rect 5000 11218 5028 12135
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5170 11112 5226 11121
rect 5170 11047 5226 11056
rect 5184 10062 5212 11047
rect 5276 10713 5304 13330
rect 5448 12844 5500 12850
rect 5552 12832 5580 14214
rect 5500 12804 5580 12832
rect 5448 12786 5500 12792
rect 5262 10704 5318 10713
rect 5262 10639 5318 10648
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5368 10577 5396 10610
rect 5354 10568 5410 10577
rect 5354 10503 5410 10512
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5368 9761 5396 10406
rect 5354 9752 5410 9761
rect 4896 9716 4948 9722
rect 5354 9687 5410 9696
rect 4896 9658 4948 9664
rect 5460 9625 5488 12786
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5446 9616 5502 9625
rect 5172 9580 5224 9586
rect 5446 9551 5502 9560
rect 5172 9522 5224 9528
rect 4724 9030 4844 9058
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4724 3534 4752 9030
rect 4986 7304 5042 7313
rect 4986 7239 5042 7248
rect 4894 7168 4950 7177
rect 4894 7103 4950 7112
rect 4802 5400 4858 5409
rect 4908 5370 4936 7103
rect 4802 5335 4858 5344
rect 4896 5364 4948 5370
rect 4816 5234 4844 5335
rect 4896 5306 4948 5312
rect 4894 5264 4950 5273
rect 4804 5228 4856 5234
rect 4894 5199 4950 5208
rect 4804 5170 4856 5176
rect 4908 4690 4936 5199
rect 5000 5098 5028 7239
rect 5078 5944 5134 5953
rect 5078 5879 5134 5888
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4908 3058 4936 4082
rect 4986 3904 5042 3913
rect 4986 3839 5042 3848
rect 5000 3194 5028 3839
rect 5092 3738 5120 5879
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5184 3670 5212 9522
rect 5552 9058 5580 11018
rect 5644 10810 5672 14470
rect 5722 14512 5778 14521
rect 5722 14447 5778 14456
rect 5736 14074 5764 14447
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5736 12345 5764 13330
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5722 12336 5778 12345
rect 5722 12271 5778 12280
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5630 10704 5686 10713
rect 5630 10639 5632 10648
rect 5684 10639 5686 10648
rect 5632 10610 5684 10616
rect 5460 9030 5580 9058
rect 5460 8974 5488 9030
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5630 8936 5686 8945
rect 5630 8871 5686 8880
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5262 8664 5318 8673
rect 5262 8599 5318 8608
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4068 2032 4120 2038
rect 4068 1974 4120 1980
rect 4344 2032 4396 2038
rect 4344 1974 4396 1980
rect 3976 1964 4028 1970
rect 3976 1906 4028 1912
rect 4250 1864 4306 1873
rect 4250 1799 4252 1808
rect 4304 1799 4306 1808
rect 4252 1770 4304 1776
rect 3146 1456 3202 1465
rect 3146 1391 3202 1400
rect 4448 1358 4476 2994
rect 5092 2446 5120 3402
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 4540 1601 4568 2382
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4804 1964 4856 1970
rect 4804 1906 4856 1912
rect 4526 1592 4582 1601
rect 4526 1527 4582 1536
rect 4816 1494 4844 1906
rect 4908 1562 4936 2246
rect 5092 1970 5120 2382
rect 5080 1964 5132 1970
rect 5080 1906 5132 1912
rect 4896 1556 4948 1562
rect 4896 1498 4948 1504
rect 4804 1488 4856 1494
rect 4804 1430 4856 1436
rect 5092 1358 5120 1906
rect 5276 1358 5304 8599
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5368 6390 5396 7482
rect 5552 6914 5580 8774
rect 5644 8498 5672 8871
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5460 6886 5580 6914
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5460 2106 5488 6886
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 5914 5580 6598
rect 5644 6254 5672 6734
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 5166 5580 5510
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5552 4826 5580 5102
rect 5644 5001 5672 6054
rect 5736 5953 5764 12106
rect 5828 11830 5856 12718
rect 6012 12209 6040 16200
rect 6472 15201 6500 16200
rect 13726 16144 13782 16153
rect 13726 16079 13782 16088
rect 9126 16008 9182 16017
rect 9126 15943 9182 15952
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 7566 15804 7874 15813
rect 7566 15802 7572 15804
rect 7628 15802 7652 15804
rect 7708 15802 7732 15804
rect 7788 15802 7812 15804
rect 7868 15802 7874 15804
rect 7628 15750 7630 15802
rect 7810 15750 7812 15802
rect 7566 15748 7572 15750
rect 7628 15748 7652 15750
rect 7708 15748 7732 15750
rect 7788 15748 7812 15750
rect 7868 15748 7874 15750
rect 7566 15739 7874 15748
rect 8114 15600 8170 15609
rect 8114 15535 8116 15544
rect 8168 15535 8170 15544
rect 8116 15506 8168 15512
rect 8392 15496 8444 15502
rect 6642 15464 6698 15473
rect 8392 15438 8444 15444
rect 6642 15399 6698 15408
rect 7380 15428 7432 15434
rect 6458 15192 6514 15201
rect 6458 15127 6514 15136
rect 6656 13938 6684 15399
rect 7380 15370 7432 15376
rect 8024 15428 8076 15434
rect 8024 15370 8076 15376
rect 7392 15094 7420 15370
rect 7380 15088 7432 15094
rect 7380 15030 7432 15036
rect 7012 14340 7064 14346
rect 7012 14282 7064 14288
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6368 12776 6420 12782
rect 6656 12753 6684 13194
rect 6368 12718 6420 12724
rect 6642 12744 6698 12753
rect 6380 12434 6408 12718
rect 6642 12679 6698 12688
rect 6288 12406 6408 12434
rect 6828 12436 6880 12442
rect 5998 12200 6054 12209
rect 5998 12135 6054 12144
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 6288 11694 6316 12406
rect 6932 12434 6960 13194
rect 6880 12406 6960 12434
rect 6828 12378 6880 12384
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6840 11801 6868 12174
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6826 11792 6882 11801
rect 6826 11727 6882 11736
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 5998 10160 6054 10169
rect 5998 10095 6000 10104
rect 6052 10095 6054 10104
rect 6000 10066 6052 10072
rect 5814 9616 5870 9625
rect 5814 9551 5870 9560
rect 5828 9518 5856 9551
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5998 9072 6054 9081
rect 5998 9007 6054 9016
rect 5906 7576 5962 7585
rect 5906 7511 5962 7520
rect 5814 6760 5870 6769
rect 5814 6695 5870 6704
rect 5828 6458 5856 6695
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5814 6352 5870 6361
rect 5814 6287 5870 6296
rect 5722 5944 5778 5953
rect 5722 5879 5778 5888
rect 5828 5302 5856 6287
rect 5920 6089 5948 7511
rect 5906 6080 5962 6089
rect 5906 6015 5962 6024
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5630 4992 5686 5001
rect 5630 4927 5686 4936
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5630 4448 5686 4457
rect 5630 4383 5686 4392
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3641 5580 3878
rect 5538 3632 5594 3641
rect 5538 3567 5594 3576
rect 5538 3496 5594 3505
rect 5538 3431 5594 3440
rect 5552 3058 5580 3431
rect 5644 3126 5672 4383
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5736 3058 5764 3402
rect 5920 3097 5948 3470
rect 6012 3194 6040 9007
rect 6288 8838 6316 11630
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6380 8537 6408 10542
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6472 8634 6500 9998
rect 6656 9926 6684 11630
rect 6828 10668 6880 10674
rect 6932 10656 6960 12038
rect 6880 10628 6960 10656
rect 6828 10610 6880 10616
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6828 9920 6880 9926
rect 6880 9880 6960 9908
rect 6828 9862 6880 9868
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6840 9489 6868 9522
rect 6826 9480 6882 9489
rect 6826 9415 6882 9424
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 9081 6776 9318
rect 6734 9072 6790 9081
rect 6734 9007 6790 9016
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6366 8528 6422 8537
rect 6366 8463 6422 8472
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6104 4826 6132 6734
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6196 5234 6224 5850
rect 6288 5681 6316 7686
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6380 7041 6408 7278
rect 6366 7032 6422 7041
rect 6366 6967 6422 6976
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6274 5672 6330 5681
rect 6274 5607 6330 5616
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6288 4622 6316 5607
rect 6472 5370 6500 6734
rect 6564 5409 6592 8910
rect 6748 8430 6776 9007
rect 6826 8528 6882 8537
rect 6932 8498 6960 9880
rect 7024 9654 7052 14282
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7116 13938 7144 14214
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7392 13410 7420 15030
rect 7566 14716 7874 14725
rect 7566 14714 7572 14716
rect 7628 14714 7652 14716
rect 7708 14714 7732 14716
rect 7788 14714 7812 14716
rect 7868 14714 7874 14716
rect 7628 14662 7630 14714
rect 7810 14662 7812 14714
rect 7566 14660 7572 14662
rect 7628 14660 7652 14662
rect 7708 14660 7732 14662
rect 7788 14660 7812 14662
rect 7868 14660 7874 14662
rect 7566 14651 7874 14660
rect 7566 13628 7874 13637
rect 7566 13626 7572 13628
rect 7628 13626 7652 13628
rect 7708 13626 7732 13628
rect 7788 13626 7812 13628
rect 7868 13626 7874 13628
rect 7628 13574 7630 13626
rect 7810 13574 7812 13626
rect 7566 13572 7572 13574
rect 7628 13572 7652 13574
rect 7708 13572 7732 13574
rect 7788 13572 7812 13574
rect 7868 13572 7874 13574
rect 7566 13563 7874 13572
rect 8036 13530 8064 15370
rect 8404 15337 8432 15438
rect 8390 15328 8446 15337
rect 8390 15263 8446 15272
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 8114 14920 8170 14929
rect 8114 14855 8170 14864
rect 8128 14521 8156 14855
rect 8114 14512 8170 14521
rect 8114 14447 8170 14456
rect 8220 14414 8248 15030
rect 8392 14952 8444 14958
rect 8390 14920 8392 14929
rect 8444 14920 8446 14929
rect 8390 14855 8446 14864
rect 8208 14408 8260 14414
rect 8260 14356 8340 14362
rect 8208 14350 8340 14356
rect 8220 14334 8340 14350
rect 8116 14000 8168 14006
rect 8114 13968 8116 13977
rect 8168 13968 8170 13977
rect 8114 13903 8170 13912
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 7300 13382 7420 13410
rect 7930 13424 7986 13433
rect 7300 12918 7328 13382
rect 7930 13359 7986 13368
rect 7944 13326 7972 13359
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 7288 12912 7340 12918
rect 8220 12889 8248 13126
rect 8312 12986 8340 14334
rect 8392 14340 8444 14346
rect 8392 14282 8444 14288
rect 8404 14249 8432 14282
rect 8390 14240 8446 14249
rect 8390 14175 8446 14184
rect 8390 13832 8446 13841
rect 8390 13767 8446 13776
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 7288 12854 7340 12860
rect 8022 12880 8078 12889
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7208 12306 7236 12718
rect 7300 12646 7328 12854
rect 8022 12815 8078 12824
rect 8206 12880 8262 12889
rect 8206 12815 8262 12824
rect 7288 12640 7340 12646
rect 7286 12608 7288 12617
rect 7932 12640 7984 12646
rect 7340 12608 7342 12617
rect 8036 12617 8064 12815
rect 7932 12582 7984 12588
rect 8022 12608 8078 12617
rect 7286 12543 7342 12552
rect 7300 12517 7328 12543
rect 7566 12540 7874 12549
rect 7566 12538 7572 12540
rect 7628 12538 7652 12540
rect 7708 12538 7732 12540
rect 7788 12538 7812 12540
rect 7868 12538 7874 12540
rect 7628 12486 7630 12538
rect 7810 12486 7812 12538
rect 7566 12484 7572 12486
rect 7628 12484 7652 12486
rect 7708 12484 7732 12486
rect 7788 12484 7812 12486
rect 7868 12484 7874 12486
rect 7566 12475 7874 12484
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7944 11898 7972 12582
rect 8022 12543 8078 12552
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8128 11898 8156 12242
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7116 11121 7144 11766
rect 7194 11656 7250 11665
rect 7194 11591 7250 11600
rect 7208 11150 7236 11591
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 7566 11452 7874 11461
rect 7566 11450 7572 11452
rect 7628 11450 7652 11452
rect 7708 11450 7732 11452
rect 7788 11450 7812 11452
rect 7868 11450 7874 11452
rect 7628 11398 7630 11450
rect 7810 11398 7812 11450
rect 7566 11396 7572 11398
rect 7628 11396 7652 11398
rect 7708 11396 7732 11398
rect 7788 11396 7812 11398
rect 7868 11396 7874 11398
rect 7566 11387 7874 11396
rect 8208 11280 8260 11286
rect 8206 11248 8208 11257
rect 8260 11248 8262 11257
rect 8206 11183 8262 11192
rect 7196 11144 7248 11150
rect 7102 11112 7158 11121
rect 7196 11086 7248 11092
rect 7102 11047 7158 11056
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 6826 8463 6882 8472
rect 6920 8492 6972 8498
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6840 8362 6868 8463
rect 6920 8434 6972 8440
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 7024 7886 7052 9590
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6642 6896 6698 6905
rect 6642 6831 6698 6840
rect 6550 5400 6606 5409
rect 6460 5364 6512 5370
rect 6550 5335 6606 5344
rect 6460 5306 6512 5312
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6090 4312 6146 4321
rect 6090 4247 6146 4256
rect 6104 3738 6132 4247
rect 6274 4176 6330 4185
rect 6274 4111 6330 4120
rect 6288 4010 6316 4111
rect 6564 4078 6592 5335
rect 6656 4690 6684 6831
rect 6748 5370 6776 7278
rect 7024 6322 7052 7686
rect 7116 7585 7144 9930
rect 7208 8265 7236 10678
rect 7194 8256 7250 8265
rect 7194 8191 7250 8200
rect 7102 7576 7158 7585
rect 7102 7511 7158 7520
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7116 7177 7144 7414
rect 7102 7168 7158 7177
rect 7102 7103 7158 7112
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6826 5808 6882 5817
rect 6826 5743 6828 5752
rect 6880 5743 6882 5752
rect 6828 5714 6880 5720
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6564 3602 6592 4014
rect 6748 3754 6776 5170
rect 6656 3726 6776 3754
rect 6840 3738 6868 5510
rect 6932 4826 6960 6190
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6918 4584 6974 4593
rect 6918 4519 6974 4528
rect 6828 3732 6880 3738
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6656 3534 6684 3726
rect 6828 3674 6880 3680
rect 6932 3618 6960 4519
rect 7024 4146 7052 5102
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7208 3738 7236 6666
rect 7300 6458 7328 11018
rect 8036 10538 8064 11018
rect 8208 10668 8260 10674
rect 8128 10628 8208 10656
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 7566 10364 7874 10373
rect 7566 10362 7572 10364
rect 7628 10362 7652 10364
rect 7708 10362 7732 10364
rect 7788 10362 7812 10364
rect 7868 10362 7874 10364
rect 7628 10310 7630 10362
rect 7810 10310 7812 10362
rect 7566 10308 7572 10310
rect 7628 10308 7652 10310
rect 7708 10308 7732 10310
rect 7788 10308 7812 10310
rect 7868 10308 7874 10310
rect 7566 10299 7874 10308
rect 8022 10024 8078 10033
rect 8022 9959 8078 9968
rect 8036 9926 8064 9959
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7566 9276 7874 9285
rect 7566 9274 7572 9276
rect 7628 9274 7652 9276
rect 7708 9274 7732 9276
rect 7788 9274 7812 9276
rect 7868 9274 7874 9276
rect 7628 9222 7630 9274
rect 7810 9222 7812 9274
rect 7566 9220 7572 9222
rect 7628 9220 7652 9222
rect 7708 9220 7732 9222
rect 7788 9220 7812 9222
rect 7868 9220 7874 9222
rect 7566 9211 7874 9220
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7392 7313 7420 8842
rect 7566 8188 7874 8197
rect 7566 8186 7572 8188
rect 7628 8186 7652 8188
rect 7708 8186 7732 8188
rect 7788 8186 7812 8188
rect 7868 8186 7874 8188
rect 7628 8134 7630 8186
rect 7810 8134 7812 8186
rect 7566 8132 7572 8134
rect 7628 8132 7652 8134
rect 7708 8132 7732 8134
rect 7788 8132 7812 8134
rect 7868 8132 7874 8134
rect 7566 8123 7874 8132
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8036 7546 8064 7822
rect 8128 7562 8156 10628
rect 8208 10610 8260 10616
rect 8206 9208 8262 9217
rect 8206 9143 8262 9152
rect 8220 8430 8248 9143
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8312 7721 8340 11494
rect 8404 9926 8432 13767
rect 8496 13569 8524 15846
rect 9140 15706 9168 15943
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 8566 15260 8874 15269
rect 8566 15258 8572 15260
rect 8628 15258 8652 15260
rect 8708 15258 8732 15260
rect 8788 15258 8812 15260
rect 8868 15258 8874 15260
rect 8628 15206 8630 15258
rect 8810 15206 8812 15258
rect 8566 15204 8572 15206
rect 8628 15204 8652 15206
rect 8708 15204 8732 15206
rect 8788 15204 8812 15206
rect 8868 15204 8874 15206
rect 8566 15195 8874 15204
rect 13358 15056 13414 15065
rect 9864 15020 9916 15026
rect 13358 14991 13414 15000
rect 9864 14962 9916 14968
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9232 14657 9260 14758
rect 9218 14648 9274 14657
rect 9218 14583 9274 14592
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 8566 14172 8874 14181
rect 8566 14170 8572 14172
rect 8628 14170 8652 14172
rect 8708 14170 8732 14172
rect 8788 14170 8812 14172
rect 8868 14170 8874 14172
rect 8628 14118 8630 14170
rect 8810 14118 8812 14170
rect 8566 14116 8572 14118
rect 8628 14116 8652 14118
rect 8708 14116 8732 14118
rect 8788 14116 8812 14118
rect 8868 14116 8874 14118
rect 8566 14107 8874 14116
rect 9232 14074 9260 14282
rect 9312 14272 9364 14278
rect 9310 14240 9312 14249
rect 9364 14240 9366 14249
rect 9310 14175 9366 14184
rect 9586 14104 9642 14113
rect 9220 14068 9272 14074
rect 9586 14039 9642 14048
rect 9220 14010 9272 14016
rect 8944 13864 8996 13870
rect 8942 13832 8944 13841
rect 8996 13832 8998 13841
rect 8942 13767 8998 13776
rect 8942 13696 8998 13705
rect 8942 13631 8998 13640
rect 8482 13560 8538 13569
rect 8482 13495 8538 13504
rect 8956 13326 8984 13631
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 9126 13288 9182 13297
rect 9126 13223 9182 13232
rect 9140 13190 9168 13223
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 8566 13084 8874 13093
rect 8566 13082 8572 13084
rect 8628 13082 8652 13084
rect 8708 13082 8732 13084
rect 8788 13082 8812 13084
rect 8868 13082 8874 13084
rect 8628 13030 8630 13082
rect 8810 13030 8812 13082
rect 8566 13028 8572 13030
rect 8628 13028 8652 13030
rect 8708 13028 8732 13030
rect 8788 13028 8812 13030
rect 8868 13028 8874 13030
rect 8566 13019 8874 13028
rect 9034 13016 9090 13025
rect 9232 13002 9260 14010
rect 9600 13938 9628 14039
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9034 12951 9090 12960
rect 9140 12974 9260 13002
rect 9048 12730 9076 12951
rect 8956 12702 9076 12730
rect 8956 12481 8984 12702
rect 9140 12594 9168 12974
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9048 12566 9168 12594
rect 8942 12472 8998 12481
rect 8942 12407 8998 12416
rect 9048 12238 9076 12566
rect 9232 12481 9260 12786
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9218 12472 9274 12481
rect 9128 12436 9180 12442
rect 9218 12407 9274 12416
rect 9128 12378 9180 12384
rect 8944 12232 8996 12238
rect 8942 12200 8944 12209
rect 9036 12232 9088 12238
rect 8996 12200 8998 12209
rect 9036 12174 9088 12180
rect 8942 12135 8998 12144
rect 8566 11996 8874 12005
rect 8566 11994 8572 11996
rect 8628 11994 8652 11996
rect 8708 11994 8732 11996
rect 8788 11994 8812 11996
rect 8868 11994 8874 11996
rect 8628 11942 8630 11994
rect 8810 11942 8812 11994
rect 8566 11940 8572 11942
rect 8628 11940 8652 11942
rect 8708 11940 8732 11942
rect 8788 11940 8812 11942
rect 8868 11940 8874 11942
rect 8566 11931 8874 11940
rect 9140 11898 9168 12378
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8390 9752 8446 9761
rect 8390 9687 8446 9696
rect 8298 7712 8354 7721
rect 8298 7647 8354 7656
rect 8128 7546 8340 7562
rect 8024 7540 8076 7546
rect 8128 7540 8352 7546
rect 8128 7534 8300 7540
rect 8024 7482 8076 7488
rect 8300 7482 8352 7488
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7378 7304 7434 7313
rect 7378 7239 7434 7248
rect 7566 7100 7874 7109
rect 7566 7098 7572 7100
rect 7628 7098 7652 7100
rect 7708 7098 7732 7100
rect 7788 7098 7812 7100
rect 7868 7098 7874 7100
rect 7628 7046 7630 7098
rect 7810 7046 7812 7098
rect 7566 7044 7572 7046
rect 7628 7044 7652 7046
rect 7708 7044 7732 7046
rect 7788 7044 7812 7046
rect 7868 7044 7874 7046
rect 7566 7035 7874 7044
rect 8036 6882 8064 7346
rect 8300 6928 8352 6934
rect 7944 6854 8064 6882
rect 8128 6876 8300 6882
rect 8128 6870 8352 6876
rect 8128 6854 8340 6870
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7286 5808 7342 5817
rect 7286 5743 7342 5752
rect 7300 5302 7328 5743
rect 7392 5574 7420 6326
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 6748 3590 6960 3618
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6748 3194 6776 3590
rect 6918 3496 6974 3505
rect 6918 3431 6974 3440
rect 6932 3194 6960 3431
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 5906 3088 5962 3097
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5724 3052 5776 3058
rect 5906 3023 5962 3032
rect 5724 2994 5776 3000
rect 7300 2825 7328 3878
rect 7286 2816 7342 2825
rect 7286 2751 7342 2760
rect 6918 2544 6974 2553
rect 7392 2514 7420 5238
rect 7484 5234 7512 6394
rect 7566 6012 7874 6021
rect 7566 6010 7572 6012
rect 7628 6010 7652 6012
rect 7708 6010 7732 6012
rect 7788 6010 7812 6012
rect 7868 6010 7874 6012
rect 7628 5958 7630 6010
rect 7810 5958 7812 6010
rect 7566 5956 7572 5958
rect 7628 5956 7652 5958
rect 7708 5956 7732 5958
rect 7788 5956 7812 5958
rect 7868 5956 7874 5958
rect 7566 5947 7874 5956
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 3058 7512 4966
rect 7566 4924 7874 4933
rect 7566 4922 7572 4924
rect 7628 4922 7652 4924
rect 7708 4922 7732 4924
rect 7788 4922 7812 4924
rect 7868 4922 7874 4924
rect 7628 4870 7630 4922
rect 7810 4870 7812 4922
rect 7566 4868 7572 4870
rect 7628 4868 7652 4870
rect 7708 4868 7732 4870
rect 7788 4868 7812 4870
rect 7868 4868 7874 4870
rect 7566 4859 7874 4868
rect 7944 4185 7972 6854
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 7930 4176 7986 4185
rect 7930 4111 7986 4120
rect 7566 3836 7874 3845
rect 7566 3834 7572 3836
rect 7628 3834 7652 3836
rect 7708 3834 7732 3836
rect 7788 3834 7812 3836
rect 7868 3834 7874 3836
rect 7628 3782 7630 3834
rect 7810 3782 7812 3834
rect 7566 3780 7572 3782
rect 7628 3780 7652 3782
rect 7708 3780 7732 3782
rect 7788 3780 7812 3782
rect 7868 3780 7874 3782
rect 7566 3771 7874 3780
rect 8036 3738 8064 6734
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8128 3534 8156 6854
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8206 5944 8262 5953
rect 8206 5879 8262 5888
rect 8220 5778 8248 5879
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8206 5672 8262 5681
rect 8206 5607 8208 5616
rect 8260 5607 8262 5616
rect 8208 5578 8260 5584
rect 8312 5114 8340 6734
rect 8404 5710 8432 9687
rect 8496 9625 8524 11086
rect 8566 10908 8874 10917
rect 8566 10906 8572 10908
rect 8628 10906 8652 10908
rect 8708 10906 8732 10908
rect 8788 10906 8812 10908
rect 8868 10906 8874 10908
rect 8628 10854 8630 10906
rect 8810 10854 8812 10906
rect 8566 10852 8572 10854
rect 8628 10852 8652 10854
rect 8708 10852 8732 10854
rect 8788 10852 8812 10854
rect 8868 10852 8874 10854
rect 8566 10843 8874 10852
rect 8956 10266 8984 11698
rect 9232 11393 9260 11698
rect 9034 11384 9090 11393
rect 9034 11319 9090 11328
rect 9218 11384 9274 11393
rect 9218 11319 9274 11328
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8566 9820 8874 9829
rect 8566 9818 8572 9820
rect 8628 9818 8652 9820
rect 8708 9818 8732 9820
rect 8788 9818 8812 9820
rect 8868 9818 8874 9820
rect 8628 9766 8630 9818
rect 8810 9766 8812 9818
rect 8566 9764 8572 9766
rect 8628 9764 8652 9766
rect 8708 9764 8732 9766
rect 8788 9764 8812 9766
rect 8868 9764 8874 9766
rect 8566 9755 8874 9764
rect 8482 9616 8538 9625
rect 9048 9602 9076 11319
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 9140 11121 9168 11222
rect 9126 11112 9182 11121
rect 9126 11047 9182 11056
rect 9600 11064 9628 12582
rect 9876 12434 9904 14962
rect 10138 14648 10194 14657
rect 10138 14583 10194 14592
rect 9954 13696 10010 13705
rect 9954 13631 10010 13640
rect 9968 12782 9996 13631
rect 10152 13326 10180 14583
rect 13372 14521 13400 14991
rect 13634 14784 13690 14793
rect 13634 14719 13690 14728
rect 11610 14512 11666 14521
rect 11610 14447 11666 14456
rect 13358 14512 13414 14521
rect 13358 14447 13414 14456
rect 10506 14376 10562 14385
rect 10506 14311 10562 14320
rect 10322 13968 10378 13977
rect 10322 13903 10378 13912
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10336 12986 10364 13903
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9876 12406 9996 12434
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9600 11036 9720 11064
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9128 10464 9180 10470
rect 9232 10441 9260 10950
rect 9128 10406 9180 10412
rect 9218 10432 9274 10441
rect 9140 10062 9168 10406
rect 9218 10367 9274 10376
rect 9232 10266 9260 10367
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9128 9648 9180 9654
rect 8482 9551 8538 9560
rect 8956 9574 9076 9602
rect 9126 9616 9128 9625
rect 9180 9616 9182 9625
rect 8566 8732 8874 8741
rect 8566 8730 8572 8732
rect 8628 8730 8652 8732
rect 8708 8730 8732 8732
rect 8788 8730 8812 8732
rect 8868 8730 8874 8732
rect 8628 8678 8630 8730
rect 8810 8678 8812 8730
rect 8566 8676 8572 8678
rect 8628 8676 8652 8678
rect 8708 8676 8732 8678
rect 8788 8676 8812 8678
rect 8868 8676 8874 8678
rect 8566 8667 8874 8676
rect 8956 7886 8984 9574
rect 9126 9551 9182 9560
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 8974 9076 9318
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9140 8566 9168 8774
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8566 7644 8874 7653
rect 8566 7642 8572 7644
rect 8628 7642 8652 7644
rect 8708 7642 8732 7644
rect 8788 7642 8812 7644
rect 8868 7642 8874 7644
rect 8628 7590 8630 7642
rect 8810 7590 8812 7642
rect 8566 7588 8572 7590
rect 8628 7588 8652 7590
rect 8708 7588 8732 7590
rect 8788 7588 8812 7590
rect 8868 7588 8874 7590
rect 8566 7579 8874 7588
rect 8956 6934 8984 7822
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 9140 6730 9168 7754
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 8566 6556 8874 6565
rect 8566 6554 8572 6556
rect 8628 6554 8652 6556
rect 8708 6554 8732 6556
rect 8788 6554 8812 6556
rect 8868 6554 8874 6556
rect 8628 6502 8630 6554
rect 8810 6502 8812 6554
rect 8566 6500 8572 6502
rect 8628 6500 8652 6502
rect 8708 6500 8732 6502
rect 8788 6500 8812 6502
rect 8868 6500 8874 6502
rect 8566 6491 8874 6500
rect 8956 6361 8984 6666
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 8942 6352 8998 6361
rect 8484 6316 8536 6322
rect 8942 6287 8998 6296
rect 8484 6258 8536 6264
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8220 5086 8340 5114
rect 8220 4282 8248 5086
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8220 3913 8248 4082
rect 8206 3904 8262 3913
rect 8206 3839 8262 3848
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 8114 2952 8170 2961
rect 8114 2887 8170 2896
rect 7566 2748 7874 2757
rect 7566 2746 7572 2748
rect 7628 2746 7652 2748
rect 7708 2746 7732 2748
rect 7788 2746 7812 2748
rect 7868 2746 7874 2748
rect 7628 2694 7630 2746
rect 7810 2694 7812 2746
rect 7566 2692 7572 2694
rect 7628 2692 7652 2694
rect 7708 2692 7732 2694
rect 7788 2692 7812 2694
rect 7868 2692 7874 2694
rect 7566 2683 7874 2692
rect 8022 2680 8078 2689
rect 8022 2615 8024 2624
rect 8076 2615 8078 2624
rect 8024 2586 8076 2592
rect 6918 2479 6974 2488
rect 7380 2508 7432 2514
rect 6736 2440 6788 2446
rect 6734 2408 6736 2417
rect 6788 2408 6790 2417
rect 6734 2343 6790 2352
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 5630 2136 5686 2145
rect 5448 2100 5500 2106
rect 5630 2071 5632 2080
rect 5448 2042 5500 2048
rect 5684 2071 5686 2080
rect 5632 2042 5684 2048
rect 6012 2038 6040 2246
rect 6000 2032 6052 2038
rect 6000 1974 6052 1980
rect 6090 2000 6146 2009
rect 5448 1964 5500 1970
rect 6932 1970 6960 2479
rect 7380 2450 7432 2456
rect 8128 2310 8156 2887
rect 8312 2774 8340 4966
rect 8390 4856 8446 4865
rect 8390 4791 8392 4800
rect 8444 4791 8446 4800
rect 8392 4762 8444 4768
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8404 4457 8432 4626
rect 8390 4448 8446 4457
rect 8390 4383 8446 4392
rect 8496 3194 8524 6258
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8566 5468 8874 5477
rect 8566 5466 8572 5468
rect 8628 5466 8652 5468
rect 8708 5466 8732 5468
rect 8788 5466 8812 5468
rect 8868 5466 8874 5468
rect 8628 5414 8630 5466
rect 8810 5414 8812 5466
rect 8566 5412 8572 5414
rect 8628 5412 8652 5414
rect 8708 5412 8732 5414
rect 8788 5412 8812 5414
rect 8868 5412 8874 5414
rect 8566 5403 8874 5412
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8588 4729 8616 5170
rect 8574 4720 8630 4729
rect 8574 4655 8630 4664
rect 8956 4622 8984 6054
rect 9048 5386 9076 6598
rect 9140 6458 9168 6666
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9126 6352 9182 6361
rect 9126 6287 9182 6296
rect 9140 5914 9168 6287
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9048 5358 9168 5386
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8566 4380 8874 4389
rect 8566 4378 8572 4380
rect 8628 4378 8652 4380
rect 8708 4378 8732 4380
rect 8788 4378 8812 4380
rect 8868 4378 8874 4380
rect 8628 4326 8630 4378
rect 8810 4326 8812 4378
rect 8566 4324 8572 4326
rect 8628 4324 8652 4326
rect 8708 4324 8732 4326
rect 8788 4324 8812 4326
rect 8868 4324 8874 4326
rect 8566 4315 8874 4324
rect 8566 3292 8874 3301
rect 8566 3290 8572 3292
rect 8628 3290 8652 3292
rect 8708 3290 8732 3292
rect 8788 3290 8812 3292
rect 8868 3290 8874 3292
rect 8628 3238 8630 3290
rect 8810 3238 8812 3290
rect 8566 3236 8572 3238
rect 8628 3236 8652 3238
rect 8708 3236 8732 3238
rect 8788 3236 8812 3238
rect 8868 3236 8874 3238
rect 8566 3227 8874 3236
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8220 2746 8340 2774
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 6090 1935 6092 1944
rect 5448 1906 5500 1912
rect 6144 1935 6146 1944
rect 6920 1964 6972 1970
rect 6092 1906 6144 1912
rect 6920 1906 6972 1912
rect 5460 1426 5488 1906
rect 6276 1760 6328 1766
rect 6276 1702 6328 1708
rect 6828 1760 6880 1766
rect 6828 1702 6880 1708
rect 6288 1465 6316 1702
rect 6274 1456 6330 1465
rect 5448 1420 5500 1426
rect 6840 1426 6868 1702
rect 7566 1660 7874 1669
rect 7566 1658 7572 1660
rect 7628 1658 7652 1660
rect 7708 1658 7732 1660
rect 7788 1658 7812 1660
rect 7868 1658 7874 1660
rect 7628 1606 7630 1658
rect 7810 1606 7812 1658
rect 7566 1604 7572 1606
rect 7628 1604 7652 1606
rect 7708 1604 7732 1606
rect 7788 1604 7812 1606
rect 7868 1604 7874 1606
rect 7566 1595 7874 1604
rect 6274 1391 6330 1400
rect 6828 1420 6880 1426
rect 5448 1362 5500 1368
rect 6828 1362 6880 1368
rect 8220 1358 8248 2746
rect 9048 2650 9076 5170
rect 9140 3534 9168 5358
rect 9232 4146 9260 10066
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9324 9489 9352 9930
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9310 9480 9366 9489
rect 9310 9415 9366 9424
rect 9416 8650 9444 9862
rect 9586 8800 9642 8809
rect 9586 8735 9642 8744
rect 9324 8622 9444 8650
rect 9324 5302 9352 8622
rect 9600 8430 9628 8735
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9310 4720 9366 4729
rect 9310 4655 9312 4664
rect 9364 4655 9366 4664
rect 9312 4626 9364 4632
rect 9312 4548 9364 4554
rect 9312 4490 9364 4496
rect 9324 4321 9352 4490
rect 9310 4312 9366 4321
rect 9310 4247 9366 4256
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9232 3777 9260 3878
rect 9218 3768 9274 3777
rect 9218 3703 9274 3712
rect 9416 3602 9444 7686
rect 9494 5672 9550 5681
rect 9494 5607 9550 5616
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9220 3392 9272 3398
rect 9218 3360 9220 3369
rect 9272 3360 9274 3369
rect 9218 3295 9274 3304
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9232 3097 9260 3130
rect 9218 3088 9274 3097
rect 9218 3023 9274 3032
rect 9402 2680 9458 2689
rect 9036 2644 9088 2650
rect 9402 2615 9458 2624
rect 9036 2586 9088 2592
rect 9416 2514 9444 2615
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8390 2136 8446 2145
rect 8496 2106 8524 2382
rect 8566 2204 8874 2213
rect 8566 2202 8572 2204
rect 8628 2202 8652 2204
rect 8708 2202 8732 2204
rect 8788 2202 8812 2204
rect 8868 2202 8874 2204
rect 8628 2150 8630 2202
rect 8810 2150 8812 2202
rect 8566 2148 8572 2150
rect 8628 2148 8652 2150
rect 8708 2148 8732 2150
rect 8788 2148 8812 2150
rect 8868 2148 8874 2150
rect 8566 2139 8874 2148
rect 9034 2136 9090 2145
rect 8390 2071 8446 2080
rect 8484 2100 8536 2106
rect 2964 1352 3016 1358
rect 1122 1320 1178 1329
rect 4436 1352 4488 1358
rect 2964 1294 3016 1300
rect 4250 1320 4306 1329
rect 1122 1255 1178 1264
rect 2976 1193 3004 1294
rect 4436 1294 4488 1300
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 5080 1352 5132 1358
rect 5080 1294 5132 1300
rect 5264 1352 5316 1358
rect 5264 1294 5316 1300
rect 6736 1352 6788 1358
rect 8208 1352 8260 1358
rect 6736 1294 6788 1300
rect 7378 1320 7434 1329
rect 4250 1255 4252 1264
rect 4304 1255 4306 1264
rect 4252 1226 4304 1232
rect 4068 1216 4120 1222
rect 846 1184 902 1193
rect 846 1119 902 1128
rect 2962 1184 3018 1193
rect 4068 1158 4120 1164
rect 2962 1119 3018 1128
rect 3566 1116 3874 1125
rect 3566 1114 3572 1116
rect 3628 1114 3652 1116
rect 3708 1114 3732 1116
rect 3788 1114 3812 1116
rect 3868 1114 3874 1116
rect 3628 1062 3630 1114
rect 3810 1062 3812 1114
rect 3566 1060 3572 1062
rect 3628 1060 3652 1062
rect 3708 1060 3732 1062
rect 3788 1060 3812 1062
rect 3868 1060 3874 1062
rect 3566 1051 3874 1060
rect 294 776 350 785
rect 294 711 350 720
rect 4080 377 4108 1158
rect 4816 921 4844 1294
rect 4988 1216 5040 1222
rect 4988 1158 5040 1164
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 6552 1216 6604 1222
rect 6552 1158 6604 1164
rect 4802 912 4858 921
rect 4802 847 4858 856
rect 5000 649 5028 1158
rect 4986 640 5042 649
rect 4986 575 5042 584
rect 4066 368 4122 377
rect 4066 303 4122 312
rect 6104 105 6132 1158
rect 6564 513 6592 1158
rect 6748 785 6776 1294
rect 8208 1294 8260 1300
rect 7378 1255 7434 1264
rect 7392 1222 7420 1255
rect 7380 1216 7432 1222
rect 7380 1158 7432 1164
rect 8404 785 8432 2071
rect 9508 2106 9536 5607
rect 9034 2071 9090 2080
rect 9496 2100 9548 2106
rect 8484 2042 8536 2048
rect 9048 2038 9076 2071
rect 9496 2042 9548 2048
rect 9036 2032 9088 2038
rect 9036 1974 9088 1980
rect 9600 1970 9628 8366
rect 9692 2774 9720 11036
rect 9784 7410 9812 12038
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9876 9897 9904 11018
rect 9862 9888 9918 9897
rect 9862 9823 9918 9832
rect 9968 9081 9996 12406
rect 10520 11966 10548 14311
rect 10690 14104 10746 14113
rect 10690 14039 10746 14048
rect 10508 11960 10560 11966
rect 10508 11902 10560 11908
rect 10704 11830 10732 14039
rect 11150 13832 11206 13841
rect 11150 13767 11206 13776
rect 10966 13152 11022 13161
rect 10966 13087 11022 13096
rect 10980 12434 11008 13087
rect 10980 12406 11100 12434
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 11072 10713 11100 12406
rect 11164 11354 11192 13767
rect 11334 13424 11390 13433
rect 11334 13359 11390 13368
rect 11348 12434 11376 13359
rect 11256 12406 11376 12434
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11150 11248 11206 11257
rect 11150 11183 11206 11192
rect 11058 10704 11114 10713
rect 11058 10639 11114 10648
rect 11164 9761 11192 11183
rect 11150 9752 11206 9761
rect 11150 9687 11206 9696
rect 11256 9330 11284 12406
rect 11624 12209 11652 14447
rect 11978 13560 12034 13569
rect 11978 13495 12034 13504
rect 11610 12200 11666 12209
rect 11610 12135 11666 12144
rect 11334 11792 11390 11801
rect 11334 11727 11390 11736
rect 11348 11257 11376 11727
rect 11992 11529 12020 13495
rect 12714 13288 12770 13297
rect 12714 13223 12770 13232
rect 12530 12880 12586 12889
rect 12530 12815 12586 12824
rect 11978 11520 12034 11529
rect 11978 11455 12034 11464
rect 12544 11393 12572 12815
rect 12622 11520 12678 11529
rect 12622 11455 12678 11464
rect 12346 11384 12402 11393
rect 11428 11348 11480 11354
rect 12346 11319 12402 11328
rect 12530 11384 12586 11393
rect 12530 11319 12586 11328
rect 11428 11290 11480 11296
rect 11334 11248 11390 11257
rect 11334 11183 11390 11192
rect 10980 9302 11284 9330
rect 9954 9072 10010 9081
rect 9954 9007 10010 9016
rect 9862 8256 9918 8265
rect 9862 8191 9918 8200
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9784 3058 9812 7210
rect 9876 5817 9904 8191
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10138 6488 10194 6497
rect 10138 6423 10194 6432
rect 9862 5808 9918 5817
rect 9862 5743 9918 5752
rect 10152 3097 10180 6423
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10138 3088 10194 3097
rect 9772 3052 9824 3058
rect 10138 3023 10194 3032
rect 9772 2994 9824 3000
rect 9692 2746 9996 2774
rect 9968 2446 9996 2746
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 9220 1964 9272 1970
rect 9220 1906 9272 1912
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 9232 1601 9260 1906
rect 9218 1592 9274 1601
rect 9218 1527 9274 1536
rect 8944 1488 8996 1494
rect 8942 1456 8944 1465
rect 8996 1456 8998 1465
rect 8942 1391 8998 1400
rect 9128 1216 9180 1222
rect 9126 1184 9128 1193
rect 9180 1184 9182 1193
rect 8566 1116 8874 1125
rect 9126 1119 9182 1128
rect 8566 1114 8572 1116
rect 8628 1114 8652 1116
rect 8708 1114 8732 1116
rect 8788 1114 8812 1116
rect 8868 1114 8874 1116
rect 8628 1062 8630 1114
rect 8810 1062 8812 1114
rect 8566 1060 8572 1062
rect 8628 1060 8652 1062
rect 8708 1060 8732 1062
rect 8788 1060 8812 1062
rect 8868 1060 8874 1062
rect 8566 1051 8874 1060
rect 10336 785 10364 3402
rect 10612 1737 10640 6802
rect 10980 4185 11008 9302
rect 11440 8945 11468 11290
rect 12360 9674 12388 11319
rect 12530 10704 12586 10713
rect 12530 10639 12586 10648
rect 12360 9646 12480 9674
rect 11426 8936 11482 8945
rect 11426 8871 11482 8880
rect 11336 7064 11388 7070
rect 11336 7006 11388 7012
rect 10966 4176 11022 4185
rect 10966 4111 11022 4120
rect 10598 1728 10654 1737
rect 10598 1663 10654 1672
rect 11348 1329 11376 7006
rect 11440 4729 11468 8871
rect 11794 7712 11850 7721
rect 11794 7647 11850 7656
rect 11426 4720 11482 4729
rect 11426 4655 11482 4664
rect 11808 3777 11836 7647
rect 12452 5114 12480 9646
rect 12544 8265 12572 10639
rect 12530 8256 12586 8265
rect 12530 8191 12586 8200
rect 12636 6633 12664 11455
rect 12728 10713 12756 13223
rect 13450 13016 13506 13025
rect 13450 12951 13506 12960
rect 13266 12200 13322 12209
rect 13266 12135 13322 12144
rect 12898 11248 12954 11257
rect 12898 11183 12954 11192
rect 12714 10704 12770 10713
rect 12714 10639 12770 10648
rect 12714 10024 12770 10033
rect 12714 9959 12770 9968
rect 12622 6624 12678 6633
rect 12622 6559 12678 6568
rect 12530 6080 12586 6089
rect 12530 6015 12586 6024
rect 12176 5086 12480 5114
rect 11886 4448 11942 4457
rect 11886 4383 11942 4392
rect 11794 3768 11850 3777
rect 11794 3703 11850 3712
rect 11900 1465 11928 4383
rect 12176 2145 12204 5086
rect 12346 4584 12402 4593
rect 12346 4519 12402 4528
rect 12360 4298 12388 4519
rect 12544 4298 12572 6015
rect 12360 4270 12572 4298
rect 12438 4176 12494 4185
rect 12348 4140 12400 4146
rect 12438 4111 12440 4120
rect 12348 4082 12400 4088
rect 12492 4111 12494 4120
rect 12440 4082 12492 4088
rect 12360 2961 12388 4082
rect 12728 4026 12756 9959
rect 12806 9752 12862 9761
rect 12806 9687 12862 9696
rect 12452 3998 12756 4026
rect 12452 3913 12480 3998
rect 12438 3904 12494 3913
rect 12438 3839 12494 3848
rect 12622 3904 12678 3913
rect 12622 3839 12678 3848
rect 12346 2952 12402 2961
rect 12346 2887 12402 2896
rect 12530 2952 12586 2961
rect 12530 2887 12586 2896
rect 12254 2816 12310 2825
rect 12544 2802 12572 2887
rect 12310 2774 12572 2802
rect 12254 2751 12310 2760
rect 12162 2136 12218 2145
rect 12162 2071 12218 2080
rect 11886 1456 11942 1465
rect 11886 1391 11942 1400
rect 11334 1320 11390 1329
rect 11334 1255 11390 1264
rect 6734 776 6790 785
rect 6734 711 6790 720
rect 8390 776 8446 785
rect 8390 711 8446 720
rect 10322 776 10378 785
rect 10322 711 10378 720
rect 12636 513 12664 3839
rect 12820 2825 12848 9687
rect 12912 2961 12940 11183
rect 13082 9888 13138 9897
rect 13082 9823 13138 9832
rect 13096 8401 13124 9823
rect 13082 8392 13138 8401
rect 13082 8327 13138 8336
rect 13280 6730 13308 12135
rect 13464 11665 13492 12951
rect 13450 11656 13506 11665
rect 13450 11591 13506 11600
rect 13648 10849 13676 14719
rect 13740 14249 13768 16079
rect 13818 15600 13874 15609
rect 13818 15535 13874 15544
rect 13726 14240 13782 14249
rect 13726 14175 13782 14184
rect 13832 13841 13860 15535
rect 14200 14113 14228 16487
rect 16578 16144 16634 16153
rect 16578 16079 16634 16088
rect 16394 15736 16450 15745
rect 16394 15671 16450 15680
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 14370 14512 14426 14521
rect 14370 14447 14426 14456
rect 15198 14512 15254 14521
rect 15198 14447 15254 14456
rect 14002 14104 14058 14113
rect 14002 14039 14058 14048
rect 14186 14104 14242 14113
rect 14186 14039 14242 14048
rect 13818 13832 13874 13841
rect 13818 13767 13874 13776
rect 13818 12744 13874 12753
rect 13818 12679 13874 12688
rect 13726 12608 13782 12617
rect 13726 12543 13782 12552
rect 13634 10840 13690 10849
rect 13634 10775 13690 10784
rect 13450 10568 13506 10577
rect 13450 10503 13452 10512
rect 13504 10503 13506 10512
rect 13452 10474 13504 10480
rect 13740 10062 13768 12543
rect 13832 12434 13860 12679
rect 14016 12434 14044 14039
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 13832 12406 13952 12434
rect 14016 12406 14228 12434
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13832 10169 13860 12310
rect 13924 12186 13952 12406
rect 13924 12158 14136 12186
rect 13910 10432 13966 10441
rect 13910 10367 13966 10376
rect 13818 10160 13874 10169
rect 13924 10130 13952 10367
rect 13818 10095 13874 10104
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13726 9752 13782 9761
rect 13726 9687 13782 9696
rect 13542 8936 13598 8945
rect 13542 8871 13598 8880
rect 13358 7304 13414 7313
rect 13358 7239 13414 7248
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 12990 5264 13046 5273
rect 12990 5199 13046 5208
rect 12898 2952 12954 2961
rect 12898 2887 12954 2896
rect 12806 2816 12862 2825
rect 12806 2751 12862 2760
rect 13004 1193 13032 5199
rect 13372 3369 13400 7239
rect 13450 6896 13506 6905
rect 13450 6831 13506 6840
rect 13464 6633 13492 6831
rect 13450 6624 13506 6633
rect 13450 6559 13506 6568
rect 13556 6361 13584 8871
rect 13740 8809 13768 9687
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13832 9353 13860 9454
rect 13818 9344 13874 9353
rect 13818 9279 13874 9288
rect 13818 9208 13874 9217
rect 13818 9143 13874 9152
rect 13726 8800 13782 8809
rect 13726 8735 13782 8744
rect 13726 8120 13782 8129
rect 13726 8055 13782 8064
rect 13634 6896 13690 6905
rect 13634 6831 13690 6840
rect 13542 6352 13598 6361
rect 13542 6287 13598 6296
rect 13544 5500 13596 5506
rect 13544 5442 13596 5448
rect 13358 3360 13414 3369
rect 13358 3295 13414 3304
rect 13556 3233 13584 5442
rect 13648 4865 13676 6831
rect 13740 6769 13768 8055
rect 13726 6760 13782 6769
rect 13726 6695 13782 6704
rect 13726 6352 13782 6361
rect 13832 6322 13860 9143
rect 14002 8392 14058 8401
rect 14002 8327 14058 8336
rect 13910 7576 13966 7585
rect 13910 7511 13966 7520
rect 13726 6287 13782 6296
rect 13820 6316 13872 6322
rect 13740 6089 13768 6287
rect 13820 6258 13872 6264
rect 13818 6216 13874 6225
rect 13924 6202 13952 7511
rect 13874 6174 13952 6202
rect 13818 6151 13874 6160
rect 13912 6112 13964 6118
rect 13726 6080 13782 6089
rect 13912 6054 13964 6060
rect 13726 6015 13782 6024
rect 13820 6044 13872 6050
rect 13820 5986 13872 5992
rect 13832 5681 13860 5986
rect 13818 5672 13874 5681
rect 13818 5607 13874 5616
rect 13832 5137 13860 5607
rect 13818 5128 13874 5137
rect 13818 5063 13874 5072
rect 13634 4856 13690 4865
rect 13634 4791 13690 4800
rect 13818 4856 13874 4865
rect 13924 4842 13952 6054
rect 13874 4814 13952 4842
rect 13818 4791 13874 4800
rect 13910 4720 13966 4729
rect 13910 4655 13966 4664
rect 13542 3224 13598 3233
rect 13542 3159 13598 3168
rect 13924 3126 13952 4655
rect 14016 4321 14044 8327
rect 14002 4312 14058 4321
rect 14002 4247 14058 4256
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 14108 2922 14136 12158
rect 14200 5506 14228 12406
rect 14292 12374 14320 13262
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14188 5500 14240 5506
rect 14188 5442 14240 5448
rect 14096 2916 14148 2922
rect 14096 2858 14148 2864
rect 12990 1184 13046 1193
rect 12990 1119 13046 1128
rect 6550 504 6606 513
rect 6550 439 6606 448
rect 12622 504 12678 513
rect 12622 439 12678 448
rect 14292 377 14320 10474
rect 14384 10441 14412 14447
rect 15108 10940 15160 10946
rect 15108 10882 15160 10888
rect 14370 10432 14426 10441
rect 14370 10367 14426 10376
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14384 6050 14412 10066
rect 14372 6044 14424 6050
rect 14372 5986 14424 5992
rect 15120 4729 15148 10882
rect 15212 9625 15240 14447
rect 15290 12064 15346 12073
rect 15290 11999 15346 12008
rect 15198 9616 15254 9625
rect 15198 9551 15254 9560
rect 15304 9466 15332 11999
rect 15396 11665 15424 15098
rect 15566 14920 15622 14929
rect 15566 14855 15622 14864
rect 16210 14920 16266 14929
rect 16210 14855 16266 14864
rect 15474 14104 15530 14113
rect 15474 14039 15530 14048
rect 15382 11656 15438 11665
rect 15382 11591 15438 11600
rect 15382 11248 15438 11257
rect 15382 11183 15438 11192
rect 15396 9518 15424 11183
rect 15488 10946 15516 14039
rect 15476 10940 15528 10946
rect 15476 10882 15528 10888
rect 15580 10538 15608 14855
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15658 12472 15714 12481
rect 15658 12407 15714 12416
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15566 10432 15622 10441
rect 15566 10367 15622 10376
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15212 9438 15332 9466
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15106 4720 15162 4729
rect 15106 4655 15162 4664
rect 15212 3505 15240 9438
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 3913 15332 9318
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15396 6769 15424 8910
rect 15488 7993 15516 10202
rect 15580 9382 15608 10367
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15568 9240 15620 9246
rect 15568 9182 15620 9188
rect 15580 8498 15608 9182
rect 15672 8974 15700 12407
rect 15764 9246 15792 12922
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 15934 12472 15990 12481
rect 15934 12407 15990 12416
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 15752 9240 15804 9246
rect 15752 9182 15804 9188
rect 15752 9104 15804 9110
rect 15752 9046 15804 9052
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15566 8392 15622 8401
rect 15566 8327 15622 8336
rect 15474 7984 15530 7993
rect 15474 7919 15530 7928
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15382 6760 15438 6769
rect 15382 6695 15438 6704
rect 15488 6526 15516 7822
rect 15476 6520 15528 6526
rect 15476 6462 15528 6468
rect 15580 5545 15608 8327
rect 15566 5536 15622 5545
rect 15566 5471 15622 5480
rect 15290 3904 15346 3913
rect 15290 3839 15346 3848
rect 15672 3641 15700 8774
rect 15764 5574 15792 9046
rect 15856 6866 15884 11766
rect 15948 7585 15976 12407
rect 15934 7576 15990 7585
rect 15934 7511 15990 7520
rect 16040 7070 16068 12718
rect 16132 11014 16160 13330
rect 16224 12102 16252 14855
rect 16302 13288 16358 13297
rect 16302 13223 16358 13232
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16212 11960 16264 11966
rect 16212 11902 16264 11908
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16118 10840 16174 10849
rect 16118 10775 16174 10784
rect 16028 7064 16080 7070
rect 16028 7006 16080 7012
rect 16132 6882 16160 10775
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 16040 6854 16160 6882
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15856 4185 15884 6598
rect 15842 4176 15898 4185
rect 15842 4111 15898 4120
rect 15658 3632 15714 3641
rect 15658 3567 15714 3576
rect 15198 3496 15254 3505
rect 15198 3431 15254 3440
rect 14554 2680 14610 2689
rect 14554 2615 14610 2624
rect 14462 2544 14518 2553
rect 14462 2479 14518 2488
rect 14476 1737 14504 2479
rect 14568 1873 14596 2615
rect 16040 2281 16068 6854
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 16026 2272 16082 2281
rect 16026 2207 16082 2216
rect 14554 1864 14610 1873
rect 14554 1799 14610 1808
rect 14462 1728 14518 1737
rect 14462 1663 14518 1672
rect 16132 921 16160 6666
rect 16224 6662 16252 11902
rect 16316 10146 16344 13223
rect 16408 12442 16436 15671
rect 16486 15328 16542 15337
rect 16486 15263 16542 15272
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 10946 16436 12038
rect 16396 10940 16448 10946
rect 16396 10882 16448 10888
rect 16394 10840 16450 10849
rect 16394 10775 16450 10784
rect 16408 10266 16436 10775
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16316 10118 16436 10146
rect 16500 10130 16528 15263
rect 16592 15162 16620 16079
rect 16684 15434 16712 16487
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16670 15328 16726 15337
rect 16670 15263 16726 15272
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16592 11150 16620 14962
rect 16684 13394 16712 15263
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16670 13288 16726 13297
rect 16670 13223 16726 13232
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16212 6520 16264 6526
rect 16212 6462 16264 6468
rect 16224 3466 16252 6462
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16118 912 16174 921
rect 16118 847 16174 856
rect 14278 368 14334 377
rect 14278 303 14334 312
rect 16316 105 16344 9998
rect 16408 6361 16436 10118
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16488 9852 16540 9858
rect 16488 9794 16540 9800
rect 16500 8838 16528 9794
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16488 8696 16540 8702
rect 16488 8638 16540 8644
rect 16500 8401 16528 8638
rect 16592 8634 16620 10950
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16684 8514 16712 13223
rect 16592 8498 16712 8514
rect 16580 8492 16712 8498
rect 16632 8486 16712 8492
rect 16580 8434 16632 8440
rect 16672 8424 16724 8430
rect 16486 8392 16542 8401
rect 16672 8366 16724 8372
rect 16486 8327 16542 8336
rect 16488 8288 16540 8294
rect 16488 8230 16540 8236
rect 16500 7274 16528 8230
rect 16580 8220 16632 8226
rect 16580 8162 16632 8168
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16592 7154 16620 8162
rect 16500 7126 16620 7154
rect 16394 6352 16450 6361
rect 16394 6287 16450 6296
rect 16500 5953 16528 7126
rect 16580 7064 16632 7070
rect 16580 7006 16632 7012
rect 16486 5944 16542 5953
rect 16486 5879 16542 5888
rect 16592 5794 16620 7006
rect 16684 6050 16712 8366
rect 16672 6044 16724 6050
rect 16672 5986 16724 5992
rect 16670 5944 16726 5953
rect 16670 5879 16726 5888
rect 16500 5766 16620 5794
rect 16500 4049 16528 5766
rect 16684 5658 16712 5879
rect 16592 5630 16712 5658
rect 16486 4040 16542 4049
rect 16486 3975 16542 3984
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 16408 649 16436 2858
rect 16592 1601 16620 5630
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16684 1737 16712 5510
rect 16670 1728 16726 1737
rect 16670 1663 16726 1672
rect 16672 1624 16724 1630
rect 16578 1592 16634 1601
rect 16672 1566 16724 1572
rect 16578 1527 16634 1536
rect 16684 1465 16712 1566
rect 16670 1456 16726 1465
rect 16670 1391 16726 1400
rect 16394 640 16450 649
rect 16394 575 16450 584
rect 6090 96 6146 105
rect 6090 31 6146 40
rect 16302 96 16358 105
rect 16302 31 16358 40
<< via2 >>
rect 386 15408 442 15464
rect 202 10648 258 10704
rect 662 13912 718 13968
rect 478 1536 534 1592
rect 1122 13232 1178 13288
rect 1030 1400 1086 1456
rect 1582 12960 1638 13016
rect 1490 12824 1546 12880
rect 1950 9560 2006 9616
rect 2572 15802 2628 15804
rect 2652 15802 2708 15804
rect 2732 15802 2788 15804
rect 2812 15802 2868 15804
rect 2572 15750 2618 15802
rect 2618 15750 2628 15802
rect 2652 15750 2682 15802
rect 2682 15750 2694 15802
rect 2694 15750 2708 15802
rect 2732 15750 2746 15802
rect 2746 15750 2758 15802
rect 2758 15750 2788 15802
rect 2812 15750 2822 15802
rect 2822 15750 2868 15802
rect 2572 15748 2628 15750
rect 2652 15748 2708 15750
rect 2732 15748 2788 15750
rect 2812 15748 2868 15750
rect 2572 14714 2628 14716
rect 2652 14714 2708 14716
rect 2732 14714 2788 14716
rect 2812 14714 2868 14716
rect 2572 14662 2618 14714
rect 2618 14662 2628 14714
rect 2652 14662 2682 14714
rect 2682 14662 2694 14714
rect 2694 14662 2708 14714
rect 2732 14662 2746 14714
rect 2746 14662 2758 14714
rect 2758 14662 2788 14714
rect 2812 14662 2822 14714
rect 2822 14662 2868 14714
rect 2572 14660 2628 14662
rect 2652 14660 2708 14662
rect 2732 14660 2788 14662
rect 2812 14660 2868 14662
rect 2502 13776 2558 13832
rect 2572 13626 2628 13628
rect 2652 13626 2708 13628
rect 2732 13626 2788 13628
rect 2812 13626 2868 13628
rect 2572 13574 2618 13626
rect 2618 13574 2628 13626
rect 2652 13574 2682 13626
rect 2682 13574 2694 13626
rect 2694 13574 2708 13626
rect 2732 13574 2746 13626
rect 2746 13574 2758 13626
rect 2758 13574 2788 13626
rect 2812 13574 2822 13626
rect 2822 13574 2868 13626
rect 2572 13572 2628 13574
rect 2652 13572 2708 13574
rect 2732 13572 2788 13574
rect 2812 13572 2868 13574
rect 2502 12724 2504 12744
rect 2504 12724 2556 12744
rect 2556 12724 2558 12744
rect 2502 12688 2558 12724
rect 2572 12538 2628 12540
rect 2652 12538 2708 12540
rect 2732 12538 2788 12540
rect 2812 12538 2868 12540
rect 2572 12486 2618 12538
rect 2618 12486 2628 12538
rect 2652 12486 2682 12538
rect 2682 12486 2694 12538
rect 2694 12486 2708 12538
rect 2732 12486 2746 12538
rect 2746 12486 2758 12538
rect 2758 12486 2788 12538
rect 2812 12486 2822 12538
rect 2822 12486 2868 12538
rect 2572 12484 2628 12486
rect 2652 12484 2708 12486
rect 2732 12484 2788 12486
rect 2812 12484 2868 12486
rect 2686 12280 2742 12336
rect 4066 16496 4122 16552
rect 3572 15258 3628 15260
rect 3652 15258 3708 15260
rect 3732 15258 3788 15260
rect 3812 15258 3868 15260
rect 3572 15206 3618 15258
rect 3618 15206 3628 15258
rect 3652 15206 3682 15258
rect 3682 15206 3694 15258
rect 3694 15206 3708 15258
rect 3732 15206 3746 15258
rect 3746 15206 3758 15258
rect 3758 15206 3788 15258
rect 3812 15206 3822 15258
rect 3822 15206 3868 15258
rect 3572 15204 3628 15206
rect 3652 15204 3708 15206
rect 3732 15204 3788 15206
rect 3812 15204 3868 15206
rect 3882 14320 3938 14376
rect 3572 14170 3628 14172
rect 3652 14170 3708 14172
rect 3732 14170 3788 14172
rect 3812 14170 3868 14172
rect 3572 14118 3618 14170
rect 3618 14118 3628 14170
rect 3652 14118 3682 14170
rect 3682 14118 3694 14170
rect 3694 14118 3708 14170
rect 3732 14118 3746 14170
rect 3746 14118 3758 14170
rect 3758 14118 3788 14170
rect 3812 14118 3822 14170
rect 3822 14118 3868 14170
rect 3572 14116 3628 14118
rect 3652 14116 3708 14118
rect 3732 14116 3788 14118
rect 3812 14116 3868 14118
rect 3330 13948 3332 13968
rect 3332 13948 3384 13968
rect 3384 13948 3386 13968
rect 3330 13912 3386 13948
rect 3238 13640 3294 13696
rect 3054 12960 3110 13016
rect 3238 12416 3294 12472
rect 2318 12144 2374 12200
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2226 10684 2228 10704
rect 2228 10684 2280 10704
rect 2280 10684 2282 10704
rect 2226 10648 2282 10684
rect 2410 10668 2466 10704
rect 2410 10648 2412 10668
rect 2412 10648 2464 10668
rect 2464 10648 2466 10668
rect 1766 8356 1822 8392
rect 1766 8336 1768 8356
rect 1768 8336 1820 8356
rect 1820 8336 1822 8356
rect 1490 6180 1546 6216
rect 1490 6160 1492 6180
rect 1492 6160 1544 6180
rect 1544 6160 1546 6180
rect 1674 4664 1730 4720
rect 2134 7792 2190 7848
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 3572 13082 3628 13084
rect 3652 13082 3708 13084
rect 3732 13082 3788 13084
rect 3812 13082 3868 13084
rect 3572 13030 3618 13082
rect 3618 13030 3628 13082
rect 3652 13030 3682 13082
rect 3682 13030 3694 13082
rect 3694 13030 3708 13082
rect 3732 13030 3746 13082
rect 3746 13030 3758 13082
rect 3758 13030 3788 13082
rect 3812 13030 3822 13082
rect 3822 13030 3868 13082
rect 3572 13028 3628 13030
rect 3652 13028 3708 13030
rect 3732 13028 3788 13030
rect 3812 13028 3868 13030
rect 3422 12824 3478 12880
rect 3882 12860 3884 12880
rect 3884 12860 3936 12880
rect 3936 12860 3938 12880
rect 3882 12824 3938 12860
rect 4158 15272 4214 15328
rect 4066 15136 4122 15192
rect 4434 15000 4490 15056
rect 4342 14900 4344 14920
rect 4344 14900 4396 14920
rect 4396 14900 4398 14920
rect 4342 14864 4398 14900
rect 4250 14184 4306 14240
rect 14186 16496 14242 16552
rect 16670 16496 16726 16552
rect 4618 15428 4674 15464
rect 4618 15408 4620 15428
rect 4620 15408 4672 15428
rect 4672 15408 4674 15428
rect 5446 16088 5502 16144
rect 5078 14184 5134 14240
rect 4894 13812 4896 13832
rect 4896 13812 4948 13832
rect 4948 13812 4950 13832
rect 4894 13776 4950 13812
rect 4526 13368 4582 13424
rect 4066 12416 4122 12472
rect 4066 12280 4122 12336
rect 3974 12008 4030 12064
rect 3572 11994 3628 11996
rect 3652 11994 3708 11996
rect 3732 11994 3788 11996
rect 3812 11994 3868 11996
rect 3572 11942 3618 11994
rect 3618 11942 3628 11994
rect 3652 11942 3682 11994
rect 3682 11942 3694 11994
rect 3694 11942 3708 11994
rect 3732 11942 3746 11994
rect 3746 11942 3758 11994
rect 3758 11942 3788 11994
rect 3812 11942 3822 11994
rect 3822 11942 3868 11994
rect 3572 11940 3628 11942
rect 3652 11940 3708 11942
rect 3732 11940 3788 11942
rect 3812 11940 3868 11942
rect 3572 10906 3628 10908
rect 3652 10906 3708 10908
rect 3732 10906 3788 10908
rect 3812 10906 3868 10908
rect 3572 10854 3618 10906
rect 3618 10854 3628 10906
rect 3652 10854 3682 10906
rect 3682 10854 3694 10906
rect 3694 10854 3708 10906
rect 3732 10854 3746 10906
rect 3746 10854 3758 10906
rect 3758 10854 3788 10906
rect 3812 10854 3822 10906
rect 3822 10854 3868 10906
rect 3572 10852 3628 10854
rect 3652 10852 3708 10854
rect 3732 10852 3788 10854
rect 3812 10852 3868 10854
rect 4342 12416 4398 12472
rect 5170 13268 5172 13288
rect 5172 13268 5224 13288
rect 5224 13268 5226 13288
rect 5170 13232 5226 13268
rect 4342 12144 4398 12200
rect 4158 11192 4214 11248
rect 4066 10104 4122 10160
rect 3572 9818 3628 9820
rect 3652 9818 3708 9820
rect 3732 9818 3788 9820
rect 3812 9818 3868 9820
rect 3572 9766 3618 9818
rect 3618 9766 3628 9818
rect 3652 9766 3682 9818
rect 3682 9766 3694 9818
rect 3694 9766 3708 9818
rect 3732 9766 3746 9818
rect 3746 9766 3758 9818
rect 3758 9766 3788 9818
rect 3812 9766 3822 9818
rect 3822 9766 3868 9818
rect 3572 9764 3628 9766
rect 3652 9764 3708 9766
rect 3732 9764 3788 9766
rect 3812 9764 3868 9766
rect 3146 8472 3202 8528
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 2226 6452 2282 6488
rect 2226 6432 2228 6452
rect 2228 6432 2280 6452
rect 2280 6432 2282 6452
rect 2226 5772 2282 5808
rect 2226 5752 2228 5772
rect 2228 5752 2280 5772
rect 2280 5752 2282 5772
rect 2962 6976 3018 7032
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 2594 5616 2650 5672
rect 2502 3984 2558 4040
rect 2410 3848 2466 3904
rect 2594 3712 2650 3768
rect 2410 3032 2466 3088
rect 2778 3712 2834 3768
rect 3572 8730 3628 8732
rect 3652 8730 3708 8732
rect 3732 8730 3788 8732
rect 3812 8730 3868 8732
rect 3572 8678 3618 8730
rect 3618 8678 3628 8730
rect 3652 8678 3682 8730
rect 3682 8678 3694 8730
rect 3694 8678 3708 8730
rect 3732 8678 3746 8730
rect 3746 8678 3758 8730
rect 3758 8678 3788 8730
rect 3812 8678 3822 8730
rect 3822 8678 3868 8730
rect 3572 8676 3628 8678
rect 3652 8676 3708 8678
rect 3732 8676 3788 8678
rect 3812 8676 3868 8678
rect 3974 8608 4030 8664
rect 3422 8336 3478 8392
rect 3238 5888 3294 5944
rect 3146 4528 3202 4584
rect 3054 4120 3110 4176
rect 2870 3440 2926 3496
rect 3330 4664 3386 4720
rect 3572 7642 3628 7644
rect 3652 7642 3708 7644
rect 3732 7642 3788 7644
rect 3812 7642 3868 7644
rect 3572 7590 3618 7642
rect 3618 7590 3628 7642
rect 3652 7590 3682 7642
rect 3682 7590 3694 7642
rect 3694 7590 3708 7642
rect 3732 7590 3746 7642
rect 3746 7590 3758 7642
rect 3758 7590 3788 7642
rect 3812 7590 3822 7642
rect 3822 7590 3868 7642
rect 3572 7588 3628 7590
rect 3652 7588 3708 7590
rect 3732 7588 3788 7590
rect 3812 7588 3868 7590
rect 3572 6554 3628 6556
rect 3652 6554 3708 6556
rect 3732 6554 3788 6556
rect 3812 6554 3868 6556
rect 3572 6502 3618 6554
rect 3618 6502 3628 6554
rect 3652 6502 3682 6554
rect 3682 6502 3694 6554
rect 3694 6502 3708 6554
rect 3732 6502 3746 6554
rect 3746 6502 3758 6554
rect 3758 6502 3788 6554
rect 3812 6502 3822 6554
rect 3822 6502 3868 6554
rect 3572 6500 3628 6502
rect 3652 6500 3708 6502
rect 3732 6500 3788 6502
rect 3812 6500 3868 6502
rect 3514 5652 3516 5672
rect 3516 5652 3568 5672
rect 3568 5652 3570 5672
rect 3514 5616 3570 5652
rect 3572 5466 3628 5468
rect 3652 5466 3708 5468
rect 3732 5466 3788 5468
rect 3812 5466 3868 5468
rect 3572 5414 3618 5466
rect 3618 5414 3628 5466
rect 3652 5414 3682 5466
rect 3682 5414 3694 5466
rect 3694 5414 3708 5466
rect 3732 5414 3746 5466
rect 3746 5414 3758 5466
rect 3758 5414 3788 5466
rect 3812 5414 3822 5466
rect 3822 5414 3868 5466
rect 3572 5412 3628 5414
rect 3652 5412 3708 5414
rect 3732 5412 3788 5414
rect 3812 5412 3868 5414
rect 3698 5072 3754 5128
rect 3572 4378 3628 4380
rect 3652 4378 3708 4380
rect 3732 4378 3788 4380
rect 3812 4378 3868 4380
rect 3572 4326 3618 4378
rect 3618 4326 3628 4378
rect 3652 4326 3682 4378
rect 3682 4326 3694 4378
rect 3694 4326 3708 4378
rect 3732 4326 3746 4378
rect 3746 4326 3758 4378
rect 3758 4326 3788 4378
rect 3812 4326 3822 4378
rect 3822 4326 3868 4378
rect 3572 4324 3628 4326
rect 3652 4324 3708 4326
rect 3732 4324 3788 4326
rect 3812 4324 3868 4326
rect 3514 3984 3570 4040
rect 3572 3290 3628 3292
rect 3652 3290 3708 3292
rect 3732 3290 3788 3292
rect 3812 3290 3868 3292
rect 3572 3238 3618 3290
rect 3618 3238 3628 3290
rect 3652 3238 3682 3290
rect 3682 3238 3694 3290
rect 3694 3238 3708 3290
rect 3732 3238 3746 3290
rect 3746 3238 3758 3290
rect 3758 3238 3788 3290
rect 3812 3238 3822 3290
rect 3822 3238 3868 3290
rect 3572 3236 3628 3238
rect 3652 3236 3708 3238
rect 3732 3236 3788 3238
rect 3812 3236 3868 3238
rect 3514 3052 3570 3088
rect 3514 3032 3516 3052
rect 3516 3032 3568 3052
rect 3568 3032 3570 3052
rect 3330 2896 3386 2952
rect 1858 1536 1914 1592
rect 2318 1536 2374 1592
rect 4158 9016 4214 9072
rect 4066 5480 4122 5536
rect 4066 4936 4122 4992
rect 4066 4020 4068 4040
rect 4068 4020 4120 4040
rect 4120 4020 4122 4040
rect 4066 3984 4122 4020
rect 4158 3712 4214 3768
rect 4526 5888 4582 5944
rect 4342 4120 4398 4176
rect 4066 2624 4122 2680
rect 3572 2202 3628 2204
rect 3652 2202 3708 2204
rect 3732 2202 3788 2204
rect 3812 2202 3868 2204
rect 3572 2150 3618 2202
rect 3618 2150 3628 2202
rect 3652 2150 3682 2202
rect 3682 2150 3694 2202
rect 3694 2150 3708 2202
rect 3732 2150 3746 2202
rect 3746 2150 3758 2202
rect 3758 2150 3788 2202
rect 3812 2150 3822 2202
rect 3822 2150 3868 2202
rect 3572 2148 3628 2150
rect 3652 2148 3708 2150
rect 3732 2148 3788 2150
rect 3812 2148 3868 2150
rect 4986 12144 5042 12200
rect 5170 11056 5226 11112
rect 5262 10648 5318 10704
rect 5354 10512 5410 10568
rect 5354 9696 5410 9752
rect 5446 9560 5502 9616
rect 4986 7248 5042 7304
rect 4894 7112 4950 7168
rect 4802 5344 4858 5400
rect 4894 5208 4950 5264
rect 5078 5888 5134 5944
rect 4986 3848 5042 3904
rect 5722 14456 5778 14512
rect 5722 12280 5778 12336
rect 5630 10668 5686 10704
rect 5630 10648 5632 10668
rect 5632 10648 5684 10668
rect 5684 10648 5686 10668
rect 5630 8880 5686 8936
rect 5262 8608 5318 8664
rect 4250 1828 4306 1864
rect 4250 1808 4252 1828
rect 4252 1808 4304 1828
rect 4304 1808 4306 1828
rect 3146 1400 3202 1456
rect 4526 1536 4582 1592
rect 13726 16088 13782 16144
rect 9126 15952 9182 16008
rect 7572 15802 7628 15804
rect 7652 15802 7708 15804
rect 7732 15802 7788 15804
rect 7812 15802 7868 15804
rect 7572 15750 7618 15802
rect 7618 15750 7628 15802
rect 7652 15750 7682 15802
rect 7682 15750 7694 15802
rect 7694 15750 7708 15802
rect 7732 15750 7746 15802
rect 7746 15750 7758 15802
rect 7758 15750 7788 15802
rect 7812 15750 7822 15802
rect 7822 15750 7868 15802
rect 7572 15748 7628 15750
rect 7652 15748 7708 15750
rect 7732 15748 7788 15750
rect 7812 15748 7868 15750
rect 8114 15564 8170 15600
rect 8114 15544 8116 15564
rect 8116 15544 8168 15564
rect 8168 15544 8170 15564
rect 6642 15408 6698 15464
rect 6458 15136 6514 15192
rect 6642 12688 6698 12744
rect 5998 12144 6054 12200
rect 6826 11736 6882 11792
rect 5998 10124 6054 10160
rect 5998 10104 6000 10124
rect 6000 10104 6052 10124
rect 6052 10104 6054 10124
rect 5814 9560 5870 9616
rect 5998 9016 6054 9072
rect 5906 7520 5962 7576
rect 5814 6704 5870 6760
rect 5814 6296 5870 6352
rect 5722 5888 5778 5944
rect 5906 6024 5962 6080
rect 5630 4936 5686 4992
rect 5630 4392 5686 4448
rect 5538 3576 5594 3632
rect 5538 3440 5594 3496
rect 6826 9424 6882 9480
rect 6734 9016 6790 9072
rect 6366 8472 6422 8528
rect 6366 6976 6422 7032
rect 6274 5616 6330 5672
rect 6826 8472 6882 8528
rect 7572 14714 7628 14716
rect 7652 14714 7708 14716
rect 7732 14714 7788 14716
rect 7812 14714 7868 14716
rect 7572 14662 7618 14714
rect 7618 14662 7628 14714
rect 7652 14662 7682 14714
rect 7682 14662 7694 14714
rect 7694 14662 7708 14714
rect 7732 14662 7746 14714
rect 7746 14662 7758 14714
rect 7758 14662 7788 14714
rect 7812 14662 7822 14714
rect 7822 14662 7868 14714
rect 7572 14660 7628 14662
rect 7652 14660 7708 14662
rect 7732 14660 7788 14662
rect 7812 14660 7868 14662
rect 7572 13626 7628 13628
rect 7652 13626 7708 13628
rect 7732 13626 7788 13628
rect 7812 13626 7868 13628
rect 7572 13574 7618 13626
rect 7618 13574 7628 13626
rect 7652 13574 7682 13626
rect 7682 13574 7694 13626
rect 7694 13574 7708 13626
rect 7732 13574 7746 13626
rect 7746 13574 7758 13626
rect 7758 13574 7788 13626
rect 7812 13574 7822 13626
rect 7822 13574 7868 13626
rect 7572 13572 7628 13574
rect 7652 13572 7708 13574
rect 7732 13572 7788 13574
rect 7812 13572 7868 13574
rect 8390 15272 8446 15328
rect 8114 14864 8170 14920
rect 8114 14456 8170 14512
rect 8390 14900 8392 14920
rect 8392 14900 8444 14920
rect 8444 14900 8446 14920
rect 8390 14864 8446 14900
rect 8114 13948 8116 13968
rect 8116 13948 8168 13968
rect 8168 13948 8170 13968
rect 8114 13912 8170 13948
rect 7930 13368 7986 13424
rect 8390 14184 8446 14240
rect 8390 13776 8446 13832
rect 8022 12824 8078 12880
rect 8206 12824 8262 12880
rect 7286 12588 7288 12608
rect 7288 12588 7340 12608
rect 7340 12588 7342 12608
rect 7286 12552 7342 12588
rect 7572 12538 7628 12540
rect 7652 12538 7708 12540
rect 7732 12538 7788 12540
rect 7812 12538 7868 12540
rect 7572 12486 7618 12538
rect 7618 12486 7628 12538
rect 7652 12486 7682 12538
rect 7682 12486 7694 12538
rect 7694 12486 7708 12538
rect 7732 12486 7746 12538
rect 7746 12486 7758 12538
rect 7758 12486 7788 12538
rect 7812 12486 7822 12538
rect 7822 12486 7868 12538
rect 7572 12484 7628 12486
rect 7652 12484 7708 12486
rect 7732 12484 7788 12486
rect 7812 12484 7868 12486
rect 8022 12552 8078 12608
rect 7194 11600 7250 11656
rect 7572 11450 7628 11452
rect 7652 11450 7708 11452
rect 7732 11450 7788 11452
rect 7812 11450 7868 11452
rect 7572 11398 7618 11450
rect 7618 11398 7628 11450
rect 7652 11398 7682 11450
rect 7682 11398 7694 11450
rect 7694 11398 7708 11450
rect 7732 11398 7746 11450
rect 7746 11398 7758 11450
rect 7758 11398 7788 11450
rect 7812 11398 7822 11450
rect 7822 11398 7868 11450
rect 7572 11396 7628 11398
rect 7652 11396 7708 11398
rect 7732 11396 7788 11398
rect 7812 11396 7868 11398
rect 8206 11228 8208 11248
rect 8208 11228 8260 11248
rect 8260 11228 8262 11248
rect 8206 11192 8262 11228
rect 7102 11056 7158 11112
rect 6642 6840 6698 6896
rect 6550 5344 6606 5400
rect 6090 4256 6146 4312
rect 6274 4120 6330 4176
rect 7194 8200 7250 8256
rect 7102 7520 7158 7576
rect 7102 7112 7158 7168
rect 6826 5772 6882 5808
rect 6826 5752 6828 5772
rect 6828 5752 6880 5772
rect 6880 5752 6882 5772
rect 6918 4528 6974 4584
rect 7572 10362 7628 10364
rect 7652 10362 7708 10364
rect 7732 10362 7788 10364
rect 7812 10362 7868 10364
rect 7572 10310 7618 10362
rect 7618 10310 7628 10362
rect 7652 10310 7682 10362
rect 7682 10310 7694 10362
rect 7694 10310 7708 10362
rect 7732 10310 7746 10362
rect 7746 10310 7758 10362
rect 7758 10310 7788 10362
rect 7812 10310 7822 10362
rect 7822 10310 7868 10362
rect 7572 10308 7628 10310
rect 7652 10308 7708 10310
rect 7732 10308 7788 10310
rect 7812 10308 7868 10310
rect 8022 9968 8078 10024
rect 7572 9274 7628 9276
rect 7652 9274 7708 9276
rect 7732 9274 7788 9276
rect 7812 9274 7868 9276
rect 7572 9222 7618 9274
rect 7618 9222 7628 9274
rect 7652 9222 7682 9274
rect 7682 9222 7694 9274
rect 7694 9222 7708 9274
rect 7732 9222 7746 9274
rect 7746 9222 7758 9274
rect 7758 9222 7788 9274
rect 7812 9222 7822 9274
rect 7822 9222 7868 9274
rect 7572 9220 7628 9222
rect 7652 9220 7708 9222
rect 7732 9220 7788 9222
rect 7812 9220 7868 9222
rect 7572 8186 7628 8188
rect 7652 8186 7708 8188
rect 7732 8186 7788 8188
rect 7812 8186 7868 8188
rect 7572 8134 7618 8186
rect 7618 8134 7628 8186
rect 7652 8134 7682 8186
rect 7682 8134 7694 8186
rect 7694 8134 7708 8186
rect 7732 8134 7746 8186
rect 7746 8134 7758 8186
rect 7758 8134 7788 8186
rect 7812 8134 7822 8186
rect 7822 8134 7868 8186
rect 7572 8132 7628 8134
rect 7652 8132 7708 8134
rect 7732 8132 7788 8134
rect 7812 8132 7868 8134
rect 8206 9152 8262 9208
rect 8572 15258 8628 15260
rect 8652 15258 8708 15260
rect 8732 15258 8788 15260
rect 8812 15258 8868 15260
rect 8572 15206 8618 15258
rect 8618 15206 8628 15258
rect 8652 15206 8682 15258
rect 8682 15206 8694 15258
rect 8694 15206 8708 15258
rect 8732 15206 8746 15258
rect 8746 15206 8758 15258
rect 8758 15206 8788 15258
rect 8812 15206 8822 15258
rect 8822 15206 8868 15258
rect 8572 15204 8628 15206
rect 8652 15204 8708 15206
rect 8732 15204 8788 15206
rect 8812 15204 8868 15206
rect 13358 15000 13414 15056
rect 9218 14592 9274 14648
rect 8572 14170 8628 14172
rect 8652 14170 8708 14172
rect 8732 14170 8788 14172
rect 8812 14170 8868 14172
rect 8572 14118 8618 14170
rect 8618 14118 8628 14170
rect 8652 14118 8682 14170
rect 8682 14118 8694 14170
rect 8694 14118 8708 14170
rect 8732 14118 8746 14170
rect 8746 14118 8758 14170
rect 8758 14118 8788 14170
rect 8812 14118 8822 14170
rect 8822 14118 8868 14170
rect 8572 14116 8628 14118
rect 8652 14116 8708 14118
rect 8732 14116 8788 14118
rect 8812 14116 8868 14118
rect 9310 14220 9312 14240
rect 9312 14220 9364 14240
rect 9364 14220 9366 14240
rect 9310 14184 9366 14220
rect 9586 14048 9642 14104
rect 8942 13812 8944 13832
rect 8944 13812 8996 13832
rect 8996 13812 8998 13832
rect 8942 13776 8998 13812
rect 8942 13640 8998 13696
rect 8482 13504 8538 13560
rect 9126 13232 9182 13288
rect 8572 13082 8628 13084
rect 8652 13082 8708 13084
rect 8732 13082 8788 13084
rect 8812 13082 8868 13084
rect 8572 13030 8618 13082
rect 8618 13030 8628 13082
rect 8652 13030 8682 13082
rect 8682 13030 8694 13082
rect 8694 13030 8708 13082
rect 8732 13030 8746 13082
rect 8746 13030 8758 13082
rect 8758 13030 8788 13082
rect 8812 13030 8822 13082
rect 8822 13030 8868 13082
rect 8572 13028 8628 13030
rect 8652 13028 8708 13030
rect 8732 13028 8788 13030
rect 8812 13028 8868 13030
rect 9034 12960 9090 13016
rect 8942 12416 8998 12472
rect 9218 12416 9274 12472
rect 8942 12180 8944 12200
rect 8944 12180 8996 12200
rect 8996 12180 8998 12200
rect 8942 12144 8998 12180
rect 8572 11994 8628 11996
rect 8652 11994 8708 11996
rect 8732 11994 8788 11996
rect 8812 11994 8868 11996
rect 8572 11942 8618 11994
rect 8618 11942 8628 11994
rect 8652 11942 8682 11994
rect 8682 11942 8694 11994
rect 8694 11942 8708 11994
rect 8732 11942 8746 11994
rect 8746 11942 8758 11994
rect 8758 11942 8788 11994
rect 8812 11942 8822 11994
rect 8822 11942 8868 11994
rect 8572 11940 8628 11942
rect 8652 11940 8708 11942
rect 8732 11940 8788 11942
rect 8812 11940 8868 11942
rect 8390 9696 8446 9752
rect 8298 7656 8354 7712
rect 7378 7248 7434 7304
rect 7572 7098 7628 7100
rect 7652 7098 7708 7100
rect 7732 7098 7788 7100
rect 7812 7098 7868 7100
rect 7572 7046 7618 7098
rect 7618 7046 7628 7098
rect 7652 7046 7682 7098
rect 7682 7046 7694 7098
rect 7694 7046 7708 7098
rect 7732 7046 7746 7098
rect 7746 7046 7758 7098
rect 7758 7046 7788 7098
rect 7812 7046 7822 7098
rect 7822 7046 7868 7098
rect 7572 7044 7628 7046
rect 7652 7044 7708 7046
rect 7732 7044 7788 7046
rect 7812 7044 7868 7046
rect 7286 5752 7342 5808
rect 6918 3440 6974 3496
rect 5906 3032 5962 3088
rect 7286 2760 7342 2816
rect 6918 2488 6974 2544
rect 7572 6010 7628 6012
rect 7652 6010 7708 6012
rect 7732 6010 7788 6012
rect 7812 6010 7868 6012
rect 7572 5958 7618 6010
rect 7618 5958 7628 6010
rect 7652 5958 7682 6010
rect 7682 5958 7694 6010
rect 7694 5958 7708 6010
rect 7732 5958 7746 6010
rect 7746 5958 7758 6010
rect 7758 5958 7788 6010
rect 7812 5958 7822 6010
rect 7822 5958 7868 6010
rect 7572 5956 7628 5958
rect 7652 5956 7708 5958
rect 7732 5956 7788 5958
rect 7812 5956 7868 5958
rect 7572 4922 7628 4924
rect 7652 4922 7708 4924
rect 7732 4922 7788 4924
rect 7812 4922 7868 4924
rect 7572 4870 7618 4922
rect 7618 4870 7628 4922
rect 7652 4870 7682 4922
rect 7682 4870 7694 4922
rect 7694 4870 7708 4922
rect 7732 4870 7746 4922
rect 7746 4870 7758 4922
rect 7758 4870 7788 4922
rect 7812 4870 7822 4922
rect 7822 4870 7868 4922
rect 7572 4868 7628 4870
rect 7652 4868 7708 4870
rect 7732 4868 7788 4870
rect 7812 4868 7868 4870
rect 7930 4120 7986 4176
rect 7572 3834 7628 3836
rect 7652 3834 7708 3836
rect 7732 3834 7788 3836
rect 7812 3834 7868 3836
rect 7572 3782 7618 3834
rect 7618 3782 7628 3834
rect 7652 3782 7682 3834
rect 7682 3782 7694 3834
rect 7694 3782 7708 3834
rect 7732 3782 7746 3834
rect 7746 3782 7758 3834
rect 7758 3782 7788 3834
rect 7812 3782 7822 3834
rect 7822 3782 7868 3834
rect 7572 3780 7628 3782
rect 7652 3780 7708 3782
rect 7732 3780 7788 3782
rect 7812 3780 7868 3782
rect 8206 5888 8262 5944
rect 8206 5636 8262 5672
rect 8206 5616 8208 5636
rect 8208 5616 8260 5636
rect 8260 5616 8262 5636
rect 8572 10906 8628 10908
rect 8652 10906 8708 10908
rect 8732 10906 8788 10908
rect 8812 10906 8868 10908
rect 8572 10854 8618 10906
rect 8618 10854 8628 10906
rect 8652 10854 8682 10906
rect 8682 10854 8694 10906
rect 8694 10854 8708 10906
rect 8732 10854 8746 10906
rect 8746 10854 8758 10906
rect 8758 10854 8788 10906
rect 8812 10854 8822 10906
rect 8822 10854 8868 10906
rect 8572 10852 8628 10854
rect 8652 10852 8708 10854
rect 8732 10852 8788 10854
rect 8812 10852 8868 10854
rect 9034 11328 9090 11384
rect 9218 11328 9274 11384
rect 8572 9818 8628 9820
rect 8652 9818 8708 9820
rect 8732 9818 8788 9820
rect 8812 9818 8868 9820
rect 8572 9766 8618 9818
rect 8618 9766 8628 9818
rect 8652 9766 8682 9818
rect 8682 9766 8694 9818
rect 8694 9766 8708 9818
rect 8732 9766 8746 9818
rect 8746 9766 8758 9818
rect 8758 9766 8788 9818
rect 8812 9766 8822 9818
rect 8822 9766 8868 9818
rect 8572 9764 8628 9766
rect 8652 9764 8708 9766
rect 8732 9764 8788 9766
rect 8812 9764 8868 9766
rect 8482 9560 8538 9616
rect 9126 11056 9182 11112
rect 10138 14592 10194 14648
rect 9954 13640 10010 13696
rect 13634 14728 13690 14784
rect 11610 14456 11666 14512
rect 13358 14456 13414 14512
rect 10506 14320 10562 14376
rect 10322 13912 10378 13968
rect 9218 10376 9274 10432
rect 9126 9596 9128 9616
rect 9128 9596 9180 9616
rect 9180 9596 9182 9616
rect 8572 8730 8628 8732
rect 8652 8730 8708 8732
rect 8732 8730 8788 8732
rect 8812 8730 8868 8732
rect 8572 8678 8618 8730
rect 8618 8678 8628 8730
rect 8652 8678 8682 8730
rect 8682 8678 8694 8730
rect 8694 8678 8708 8730
rect 8732 8678 8746 8730
rect 8746 8678 8758 8730
rect 8758 8678 8788 8730
rect 8812 8678 8822 8730
rect 8822 8678 8868 8730
rect 8572 8676 8628 8678
rect 8652 8676 8708 8678
rect 8732 8676 8788 8678
rect 8812 8676 8868 8678
rect 9126 9560 9182 9596
rect 8572 7642 8628 7644
rect 8652 7642 8708 7644
rect 8732 7642 8788 7644
rect 8812 7642 8868 7644
rect 8572 7590 8618 7642
rect 8618 7590 8628 7642
rect 8652 7590 8682 7642
rect 8682 7590 8694 7642
rect 8694 7590 8708 7642
rect 8732 7590 8746 7642
rect 8746 7590 8758 7642
rect 8758 7590 8788 7642
rect 8812 7590 8822 7642
rect 8822 7590 8868 7642
rect 8572 7588 8628 7590
rect 8652 7588 8708 7590
rect 8732 7588 8788 7590
rect 8812 7588 8868 7590
rect 8572 6554 8628 6556
rect 8652 6554 8708 6556
rect 8732 6554 8788 6556
rect 8812 6554 8868 6556
rect 8572 6502 8618 6554
rect 8618 6502 8628 6554
rect 8652 6502 8682 6554
rect 8682 6502 8694 6554
rect 8694 6502 8708 6554
rect 8732 6502 8746 6554
rect 8746 6502 8758 6554
rect 8758 6502 8788 6554
rect 8812 6502 8822 6554
rect 8822 6502 8868 6554
rect 8572 6500 8628 6502
rect 8652 6500 8708 6502
rect 8732 6500 8788 6502
rect 8812 6500 8868 6502
rect 8942 6296 8998 6352
rect 8206 3848 8262 3904
rect 8114 2896 8170 2952
rect 7572 2746 7628 2748
rect 7652 2746 7708 2748
rect 7732 2746 7788 2748
rect 7812 2746 7868 2748
rect 7572 2694 7618 2746
rect 7618 2694 7628 2746
rect 7652 2694 7682 2746
rect 7682 2694 7694 2746
rect 7694 2694 7708 2746
rect 7732 2694 7746 2746
rect 7746 2694 7758 2746
rect 7758 2694 7788 2746
rect 7812 2694 7822 2746
rect 7822 2694 7868 2746
rect 7572 2692 7628 2694
rect 7652 2692 7708 2694
rect 7732 2692 7788 2694
rect 7812 2692 7868 2694
rect 8022 2644 8078 2680
rect 8022 2624 8024 2644
rect 8024 2624 8076 2644
rect 8076 2624 8078 2644
rect 6734 2388 6736 2408
rect 6736 2388 6788 2408
rect 6788 2388 6790 2408
rect 6734 2352 6790 2388
rect 5630 2100 5686 2136
rect 5630 2080 5632 2100
rect 5632 2080 5684 2100
rect 5684 2080 5686 2100
rect 6090 1964 6146 2000
rect 8390 4820 8446 4856
rect 8390 4800 8392 4820
rect 8392 4800 8444 4820
rect 8444 4800 8446 4820
rect 8390 4392 8446 4448
rect 8572 5466 8628 5468
rect 8652 5466 8708 5468
rect 8732 5466 8788 5468
rect 8812 5466 8868 5468
rect 8572 5414 8618 5466
rect 8618 5414 8628 5466
rect 8652 5414 8682 5466
rect 8682 5414 8694 5466
rect 8694 5414 8708 5466
rect 8732 5414 8746 5466
rect 8746 5414 8758 5466
rect 8758 5414 8788 5466
rect 8812 5414 8822 5466
rect 8822 5414 8868 5466
rect 8572 5412 8628 5414
rect 8652 5412 8708 5414
rect 8732 5412 8788 5414
rect 8812 5412 8868 5414
rect 8574 4664 8630 4720
rect 9126 6296 9182 6352
rect 8572 4378 8628 4380
rect 8652 4378 8708 4380
rect 8732 4378 8788 4380
rect 8812 4378 8868 4380
rect 8572 4326 8618 4378
rect 8618 4326 8628 4378
rect 8652 4326 8682 4378
rect 8682 4326 8694 4378
rect 8694 4326 8708 4378
rect 8732 4326 8746 4378
rect 8746 4326 8758 4378
rect 8758 4326 8788 4378
rect 8812 4326 8822 4378
rect 8822 4326 8868 4378
rect 8572 4324 8628 4326
rect 8652 4324 8708 4326
rect 8732 4324 8788 4326
rect 8812 4324 8868 4326
rect 8572 3290 8628 3292
rect 8652 3290 8708 3292
rect 8732 3290 8788 3292
rect 8812 3290 8868 3292
rect 8572 3238 8618 3290
rect 8618 3238 8628 3290
rect 8652 3238 8682 3290
rect 8682 3238 8694 3290
rect 8694 3238 8708 3290
rect 8732 3238 8746 3290
rect 8746 3238 8758 3290
rect 8758 3238 8788 3290
rect 8812 3238 8822 3290
rect 8822 3238 8868 3290
rect 8572 3236 8628 3238
rect 8652 3236 8708 3238
rect 8732 3236 8788 3238
rect 8812 3236 8868 3238
rect 6090 1944 6092 1964
rect 6092 1944 6144 1964
rect 6144 1944 6146 1964
rect 6274 1400 6330 1456
rect 7572 1658 7628 1660
rect 7652 1658 7708 1660
rect 7732 1658 7788 1660
rect 7812 1658 7868 1660
rect 7572 1606 7618 1658
rect 7618 1606 7628 1658
rect 7652 1606 7682 1658
rect 7682 1606 7694 1658
rect 7694 1606 7708 1658
rect 7732 1606 7746 1658
rect 7746 1606 7758 1658
rect 7758 1606 7788 1658
rect 7812 1606 7822 1658
rect 7822 1606 7868 1658
rect 7572 1604 7628 1606
rect 7652 1604 7708 1606
rect 7732 1604 7788 1606
rect 7812 1604 7868 1606
rect 9310 9424 9366 9480
rect 9586 8744 9642 8800
rect 9310 4684 9366 4720
rect 9310 4664 9312 4684
rect 9312 4664 9364 4684
rect 9364 4664 9366 4684
rect 9310 4256 9366 4312
rect 9218 3712 9274 3768
rect 9494 5616 9550 5672
rect 9218 3340 9220 3360
rect 9220 3340 9272 3360
rect 9272 3340 9274 3360
rect 9218 3304 9274 3340
rect 9218 3032 9274 3088
rect 9402 2624 9458 2680
rect 8390 2080 8446 2136
rect 8572 2202 8628 2204
rect 8652 2202 8708 2204
rect 8732 2202 8788 2204
rect 8812 2202 8868 2204
rect 8572 2150 8618 2202
rect 8618 2150 8628 2202
rect 8652 2150 8682 2202
rect 8682 2150 8694 2202
rect 8694 2150 8708 2202
rect 8732 2150 8746 2202
rect 8746 2150 8758 2202
rect 8758 2150 8788 2202
rect 8812 2150 8822 2202
rect 8822 2150 8868 2202
rect 8572 2148 8628 2150
rect 8652 2148 8708 2150
rect 8732 2148 8788 2150
rect 8812 2148 8868 2150
rect 1122 1264 1178 1320
rect 4250 1284 4306 1320
rect 4250 1264 4252 1284
rect 4252 1264 4304 1284
rect 4304 1264 4306 1284
rect 846 1128 902 1184
rect 2962 1128 3018 1184
rect 3572 1114 3628 1116
rect 3652 1114 3708 1116
rect 3732 1114 3788 1116
rect 3812 1114 3868 1116
rect 3572 1062 3618 1114
rect 3618 1062 3628 1114
rect 3652 1062 3682 1114
rect 3682 1062 3694 1114
rect 3694 1062 3708 1114
rect 3732 1062 3746 1114
rect 3746 1062 3758 1114
rect 3758 1062 3788 1114
rect 3812 1062 3822 1114
rect 3822 1062 3868 1114
rect 3572 1060 3628 1062
rect 3652 1060 3708 1062
rect 3732 1060 3788 1062
rect 3812 1060 3868 1062
rect 294 720 350 776
rect 4802 856 4858 912
rect 4986 584 5042 640
rect 4066 312 4122 368
rect 7378 1264 7434 1320
rect 9034 2080 9090 2136
rect 9862 9832 9918 9888
rect 10690 14048 10746 14104
rect 11150 13776 11206 13832
rect 10966 13096 11022 13152
rect 11334 13368 11390 13424
rect 11150 11192 11206 11248
rect 11058 10648 11114 10704
rect 11150 9696 11206 9752
rect 11978 13504 12034 13560
rect 11610 12144 11666 12200
rect 11334 11736 11390 11792
rect 12714 13232 12770 13288
rect 12530 12824 12586 12880
rect 11978 11464 12034 11520
rect 12622 11464 12678 11520
rect 12346 11328 12402 11384
rect 12530 11328 12586 11384
rect 11334 11192 11390 11248
rect 9954 9016 10010 9072
rect 9862 8200 9918 8256
rect 10138 6432 10194 6488
rect 9862 5752 9918 5808
rect 10138 3032 10194 3088
rect 9218 1536 9274 1592
rect 8942 1436 8944 1456
rect 8944 1436 8996 1456
rect 8996 1436 8998 1456
rect 8942 1400 8998 1436
rect 9126 1164 9128 1184
rect 9128 1164 9180 1184
rect 9180 1164 9182 1184
rect 9126 1128 9182 1164
rect 8572 1114 8628 1116
rect 8652 1114 8708 1116
rect 8732 1114 8788 1116
rect 8812 1114 8868 1116
rect 8572 1062 8618 1114
rect 8618 1062 8628 1114
rect 8652 1062 8682 1114
rect 8682 1062 8694 1114
rect 8694 1062 8708 1114
rect 8732 1062 8746 1114
rect 8746 1062 8758 1114
rect 8758 1062 8788 1114
rect 8812 1062 8822 1114
rect 8822 1062 8868 1114
rect 8572 1060 8628 1062
rect 8652 1060 8708 1062
rect 8732 1060 8788 1062
rect 8812 1060 8868 1062
rect 12530 10648 12586 10704
rect 11426 8880 11482 8936
rect 10966 4120 11022 4176
rect 10598 1672 10654 1728
rect 11794 7656 11850 7712
rect 11426 4664 11482 4720
rect 12530 8200 12586 8256
rect 13450 12960 13506 13016
rect 13266 12144 13322 12200
rect 12898 11192 12954 11248
rect 12714 10648 12770 10704
rect 12714 9968 12770 10024
rect 12622 6568 12678 6624
rect 12530 6024 12586 6080
rect 11886 4392 11942 4448
rect 11794 3712 11850 3768
rect 12346 4528 12402 4584
rect 12438 4140 12494 4176
rect 12438 4120 12440 4140
rect 12440 4120 12492 4140
rect 12492 4120 12494 4140
rect 12806 9696 12862 9752
rect 12438 3848 12494 3904
rect 12622 3848 12678 3904
rect 12346 2896 12402 2952
rect 12530 2896 12586 2952
rect 12254 2760 12310 2816
rect 12162 2080 12218 2136
rect 11886 1400 11942 1456
rect 11334 1264 11390 1320
rect 6734 720 6790 776
rect 8390 720 8446 776
rect 10322 720 10378 776
rect 13082 9832 13138 9888
rect 13082 8336 13138 8392
rect 13450 11600 13506 11656
rect 13818 15544 13874 15600
rect 13726 14184 13782 14240
rect 16578 16088 16634 16144
rect 16394 15680 16450 15736
rect 14370 14456 14426 14512
rect 15198 14456 15254 14512
rect 14002 14048 14058 14104
rect 14186 14048 14242 14104
rect 13818 13776 13874 13832
rect 13818 12688 13874 12744
rect 13726 12552 13782 12608
rect 13634 10784 13690 10840
rect 13450 10532 13506 10568
rect 13450 10512 13452 10532
rect 13452 10512 13504 10532
rect 13504 10512 13506 10532
rect 13910 10376 13966 10432
rect 13818 10104 13874 10160
rect 13726 9696 13782 9752
rect 13542 8880 13598 8936
rect 13358 7248 13414 7304
rect 12990 5208 13046 5264
rect 12898 2896 12954 2952
rect 12806 2760 12862 2816
rect 13450 6840 13506 6896
rect 13450 6568 13506 6624
rect 13818 9288 13874 9344
rect 13818 9152 13874 9208
rect 13726 8744 13782 8800
rect 13726 8064 13782 8120
rect 13634 6840 13690 6896
rect 13542 6296 13598 6352
rect 13358 3304 13414 3360
rect 13726 6704 13782 6760
rect 13726 6296 13782 6352
rect 14002 8336 14058 8392
rect 13910 7520 13966 7576
rect 13818 6160 13874 6216
rect 13726 6024 13782 6080
rect 13818 5616 13874 5672
rect 13818 5072 13874 5128
rect 13634 4800 13690 4856
rect 13818 4800 13874 4856
rect 13910 4664 13966 4720
rect 13542 3168 13598 3224
rect 14002 4256 14058 4312
rect 12990 1128 13046 1184
rect 6550 448 6606 504
rect 12622 448 12678 504
rect 14370 10376 14426 10432
rect 15290 12008 15346 12064
rect 15198 9560 15254 9616
rect 15566 14864 15622 14920
rect 16210 14864 16266 14920
rect 15474 14048 15530 14104
rect 15382 11600 15438 11656
rect 15382 11192 15438 11248
rect 15658 12416 15714 12472
rect 15566 10376 15622 10432
rect 15106 4664 15162 4720
rect 15934 12416 15990 12472
rect 15566 8336 15622 8392
rect 15474 7928 15530 7984
rect 15382 6704 15438 6760
rect 15566 5480 15622 5536
rect 15290 3848 15346 3904
rect 15934 7520 15990 7576
rect 16302 13232 16358 13288
rect 16118 10784 16174 10840
rect 15842 4120 15898 4176
rect 15658 3576 15714 3632
rect 15198 3440 15254 3496
rect 14554 2624 14610 2680
rect 14462 2488 14518 2544
rect 16026 2216 16082 2272
rect 14554 1808 14610 1864
rect 14462 1672 14518 1728
rect 16486 15272 16542 15328
rect 16394 10784 16450 10840
rect 16670 15272 16726 15328
rect 16670 13232 16726 13288
rect 16118 856 16174 912
rect 14278 312 14334 368
rect 16486 8336 16542 8392
rect 16394 6296 16450 6352
rect 16486 5888 16542 5944
rect 16670 5888 16726 5944
rect 16486 3984 16542 4040
rect 16670 1672 16726 1728
rect 16578 1536 16634 1592
rect 16670 1400 16726 1456
rect 16394 584 16450 640
rect 6090 40 6146 96
rect 16302 40 16358 96
<< metal3 >>
rect 4061 16554 4127 16557
rect 14181 16554 14247 16557
rect 16665 16554 16731 16557
rect 4061 16552 14247 16554
rect 4061 16496 4066 16552
rect 4122 16496 14186 16552
rect 14242 16496 14247 16552
rect 4061 16494 14247 16496
rect 4061 16491 4127 16494
rect 14181 16491 14247 16494
rect 16622 16552 16731 16554
rect 16622 16496 16670 16552
rect 16726 16496 16731 16552
rect 16622 16491 16731 16496
rect 16622 16368 16682 16491
rect 14000 16248 34000 16368
rect 5441 16146 5507 16149
rect 13721 16146 13787 16149
rect 16573 16146 16639 16149
rect 5441 16144 13787 16146
rect 5441 16088 5446 16144
rect 5502 16088 13726 16144
rect 13782 16088 13787 16144
rect 5441 16086 13787 16088
rect 5441 16083 5507 16086
rect 13721 16083 13787 16086
rect 13862 16144 16639 16146
rect 13862 16088 16578 16144
rect 16634 16088 16639 16144
rect 13862 16086 16639 16088
rect 9121 16010 9187 16013
rect 13862 16010 13922 16086
rect 16573 16083 16639 16086
rect 9121 16008 13922 16010
rect 9121 15952 9126 16008
rect 9182 15952 13922 16008
rect 9121 15950 13922 15952
rect 9121 15947 9187 15950
rect 14000 15874 34000 15960
rect 13862 15840 34000 15874
rect 13862 15814 14076 15840
rect 2562 15808 2878 15809
rect 2562 15744 2568 15808
rect 2632 15744 2648 15808
rect 2712 15744 2728 15808
rect 2792 15744 2808 15808
rect 2872 15744 2878 15808
rect 2562 15743 2878 15744
rect 7562 15808 7878 15809
rect 7562 15744 7568 15808
rect 7632 15744 7648 15808
rect 7712 15744 7728 15808
rect 7792 15744 7808 15808
rect 7872 15744 7878 15808
rect 7562 15743 7878 15744
rect 13862 15738 13922 15814
rect 16389 15738 16455 15741
rect 13862 15736 16455 15738
rect 13862 15680 16394 15736
rect 16450 15680 16455 15736
rect 13862 15678 16455 15680
rect 16389 15675 16455 15678
rect 8109 15602 8175 15605
rect 13813 15602 13879 15605
rect 8109 15600 13879 15602
rect 8109 15544 8114 15600
rect 8170 15544 13818 15600
rect 13874 15544 13879 15600
rect 8109 15542 13879 15544
rect 8109 15539 8175 15542
rect 13813 15539 13879 15542
rect 381 15466 447 15469
rect 4613 15466 4679 15469
rect 381 15464 4679 15466
rect 381 15408 386 15464
rect 442 15408 4618 15464
rect 4674 15408 4679 15464
rect 381 15406 4679 15408
rect 381 15403 447 15406
rect 4613 15403 4679 15406
rect 6637 15466 6703 15469
rect 6637 15464 12450 15466
rect 6637 15408 6642 15464
rect 6698 15408 12450 15464
rect 14000 15432 34000 15552
rect 6637 15406 12450 15408
rect 6637 15403 6703 15406
rect 4153 15330 4219 15333
rect 8385 15330 8451 15333
rect 4153 15328 8451 15330
rect 4153 15272 4158 15328
rect 4214 15272 8390 15328
rect 8446 15272 8451 15328
rect 4153 15270 8451 15272
rect 12390 15330 12450 15406
rect 16622 15333 16682 15432
rect 16481 15330 16547 15333
rect 12390 15328 16547 15330
rect 12390 15272 16486 15328
rect 16542 15272 16547 15328
rect 12390 15270 16547 15272
rect 16622 15328 16731 15333
rect 16622 15272 16670 15328
rect 16726 15272 16731 15328
rect 16622 15270 16731 15272
rect 4153 15267 4219 15270
rect 8385 15267 8451 15270
rect 16481 15267 16547 15270
rect 16665 15267 16731 15270
rect 3562 15264 3878 15265
rect 3562 15200 3568 15264
rect 3632 15200 3648 15264
rect 3712 15200 3728 15264
rect 3792 15200 3808 15264
rect 3872 15200 3878 15264
rect 3562 15199 3878 15200
rect 8562 15264 8878 15265
rect 8562 15200 8568 15264
rect 8632 15200 8648 15264
rect 8712 15200 8728 15264
rect 8792 15200 8808 15264
rect 8872 15200 8878 15264
rect 8562 15199 8878 15200
rect 4061 15194 4127 15197
rect 6453 15194 6519 15197
rect 4061 15192 6519 15194
rect 4061 15136 4066 15192
rect 4122 15136 6458 15192
rect 6514 15136 6519 15192
rect 4061 15134 6519 15136
rect 4061 15131 4127 15134
rect 6453 15131 6519 15134
rect 4429 15058 4495 15061
rect 13353 15058 13419 15061
rect 4429 15056 13419 15058
rect 4429 15000 4434 15056
rect 4490 15000 13358 15056
rect 13414 15000 13419 15056
rect 14000 15024 34000 15144
rect 4429 14998 13419 15000
rect 4429 14995 4495 14998
rect 13353 14995 13419 14998
rect 16254 14925 16314 15024
rect 4337 14922 4403 14925
rect 8109 14922 8175 14925
rect 4337 14920 8175 14922
rect 4337 14864 4342 14920
rect 4398 14864 8114 14920
rect 8170 14864 8175 14920
rect 4337 14862 8175 14864
rect 4337 14859 4403 14862
rect 8109 14859 8175 14862
rect 8385 14922 8451 14925
rect 15561 14922 15627 14925
rect 8385 14920 15627 14922
rect 8385 14864 8390 14920
rect 8446 14864 15566 14920
rect 15622 14864 15627 14920
rect 8385 14862 15627 14864
rect 8385 14859 8451 14862
rect 15561 14859 15627 14862
rect 16205 14920 16314 14925
rect 16205 14864 16210 14920
rect 16266 14864 16314 14920
rect 16205 14862 16314 14864
rect 16205 14859 16271 14862
rect 13629 14786 13695 14789
rect 7974 14784 13695 14786
rect 7974 14728 13634 14784
rect 13690 14728 13695 14784
rect 7974 14726 13695 14728
rect 2562 14720 2878 14721
rect 2562 14656 2568 14720
rect 2632 14656 2648 14720
rect 2712 14656 2728 14720
rect 2792 14656 2808 14720
rect 2872 14656 2878 14720
rect 2562 14655 2878 14656
rect 7562 14720 7878 14721
rect 7562 14656 7568 14720
rect 7632 14656 7648 14720
rect 7712 14656 7728 14720
rect 7792 14656 7808 14720
rect 7872 14656 7878 14720
rect 7562 14655 7878 14656
rect 5717 14514 5783 14517
rect 7974 14514 8034 14726
rect 13629 14723 13695 14726
rect 9213 14650 9279 14653
rect 10133 14650 10199 14653
rect 9213 14648 10199 14650
rect 9213 14592 9218 14648
rect 9274 14592 10138 14648
rect 10194 14592 10199 14648
rect 14000 14616 34000 14736
rect 9213 14590 10199 14592
rect 9213 14587 9279 14590
rect 10133 14587 10199 14590
rect 15150 14517 15210 14616
rect 5717 14512 8034 14514
rect 5717 14456 5722 14512
rect 5778 14456 8034 14512
rect 5717 14454 8034 14456
rect 8109 14514 8175 14517
rect 11605 14514 11671 14517
rect 8109 14512 11671 14514
rect 8109 14456 8114 14512
rect 8170 14456 11610 14512
rect 11666 14456 11671 14512
rect 8109 14454 11671 14456
rect 5717 14451 5783 14454
rect 8109 14451 8175 14454
rect 11605 14451 11671 14454
rect 13353 14514 13419 14517
rect 14365 14514 14431 14517
rect 13353 14512 14431 14514
rect 13353 14456 13358 14512
rect 13414 14456 14370 14512
rect 14426 14456 14431 14512
rect 13353 14454 14431 14456
rect 15150 14512 15259 14517
rect 15150 14456 15198 14512
rect 15254 14456 15259 14512
rect 15150 14454 15259 14456
rect 13353 14451 13419 14454
rect 14365 14451 14431 14454
rect 15193 14451 15259 14454
rect 3877 14378 3943 14381
rect 10501 14378 10567 14381
rect 3877 14376 10567 14378
rect 3877 14320 3882 14376
rect 3938 14320 10506 14376
rect 10562 14320 10567 14376
rect 3877 14318 10567 14320
rect 3877 14315 3943 14318
rect 10501 14315 10567 14318
rect 4245 14242 4311 14245
rect 5073 14242 5139 14245
rect 8385 14242 8451 14245
rect 4245 14240 8451 14242
rect 4245 14184 4250 14240
rect 4306 14184 5078 14240
rect 5134 14184 8390 14240
rect 8446 14184 8451 14240
rect 4245 14182 8451 14184
rect 4245 14179 4311 14182
rect 5073 14179 5139 14182
rect 8385 14179 8451 14182
rect 9305 14242 9371 14245
rect 13721 14242 13787 14245
rect 14000 14242 34000 14328
rect 9305 14240 13186 14242
rect 9305 14184 9310 14240
rect 9366 14184 13186 14240
rect 9305 14182 13186 14184
rect 9305 14179 9371 14182
rect 3562 14176 3878 14177
rect 3562 14112 3568 14176
rect 3632 14112 3648 14176
rect 3712 14112 3728 14176
rect 3792 14112 3808 14176
rect 3872 14112 3878 14176
rect 3562 14111 3878 14112
rect 8562 14176 8878 14177
rect 8562 14112 8568 14176
rect 8632 14112 8648 14176
rect 8712 14112 8728 14176
rect 8792 14112 8808 14176
rect 8872 14112 8878 14176
rect 8562 14111 8878 14112
rect 9581 14106 9647 14109
rect 10685 14106 10751 14109
rect 9581 14104 10751 14106
rect 9581 14048 9586 14104
rect 9642 14048 10690 14104
rect 10746 14048 10751 14104
rect 9581 14046 10751 14048
rect 13126 14106 13186 14182
rect 13721 14240 34000 14242
rect 13721 14184 13726 14240
rect 13782 14208 34000 14240
rect 13782 14184 14076 14208
rect 13721 14182 14076 14184
rect 13721 14179 13787 14182
rect 13997 14106 14063 14109
rect 13126 14104 14063 14106
rect 13126 14048 14002 14104
rect 14058 14048 14063 14104
rect 13126 14046 14063 14048
rect 9581 14043 9647 14046
rect 10685 14043 10751 14046
rect 13997 14043 14063 14046
rect 14181 14106 14247 14109
rect 15469 14106 15535 14109
rect 14181 14104 15535 14106
rect 14181 14048 14186 14104
rect 14242 14048 15474 14104
rect 15530 14048 15535 14104
rect 14181 14046 15535 14048
rect 14181 14043 14247 14046
rect 15469 14043 15535 14046
rect 657 13970 723 13973
rect 3325 13970 3391 13973
rect 657 13968 3391 13970
rect 657 13912 662 13968
rect 718 13912 3330 13968
rect 3386 13912 3391 13968
rect 657 13910 3391 13912
rect 657 13907 723 13910
rect 3325 13907 3391 13910
rect 8109 13970 8175 13973
rect 10317 13970 10383 13973
rect 8109 13968 10383 13970
rect 8109 13912 8114 13968
rect 8170 13912 10322 13968
rect 10378 13912 10383 13968
rect 8109 13910 10383 13912
rect 8109 13907 8175 13910
rect 10317 13907 10383 13910
rect 2497 13834 2563 13837
rect 4889 13834 4955 13837
rect 8385 13834 8451 13837
rect 2497 13832 3250 13834
rect 2497 13776 2502 13832
rect 2558 13776 3250 13832
rect 2497 13774 3250 13776
rect 2497 13771 2563 13774
rect 3190 13701 3250 13774
rect 4889 13832 8451 13834
rect 4889 13776 4894 13832
rect 4950 13776 8390 13832
rect 8446 13776 8451 13832
rect 4889 13774 8451 13776
rect 4889 13771 4955 13774
rect 8385 13771 8451 13774
rect 8937 13834 9003 13837
rect 11145 13834 11211 13837
rect 8937 13832 11211 13834
rect 8937 13776 8942 13832
rect 8998 13776 11150 13832
rect 11206 13776 11211 13832
rect 8937 13774 11211 13776
rect 8937 13771 9003 13774
rect 11145 13771 11211 13774
rect 13813 13834 13879 13837
rect 14000 13834 34000 13920
rect 13813 13832 34000 13834
rect 13813 13776 13818 13832
rect 13874 13800 34000 13832
rect 13874 13776 14076 13800
rect 13813 13774 14076 13776
rect 13813 13771 13879 13774
rect 3190 13696 3299 13701
rect 3190 13640 3238 13696
rect 3294 13640 3299 13696
rect 3190 13638 3299 13640
rect 3233 13635 3299 13638
rect 8937 13698 9003 13701
rect 9949 13698 10015 13701
rect 8937 13696 10015 13698
rect 8937 13640 8942 13696
rect 8998 13640 9954 13696
rect 10010 13640 10015 13696
rect 8937 13638 10015 13640
rect 8937 13635 9003 13638
rect 9949 13635 10015 13638
rect 2562 13632 2878 13633
rect 2562 13568 2568 13632
rect 2632 13568 2648 13632
rect 2712 13568 2728 13632
rect 2792 13568 2808 13632
rect 2872 13568 2878 13632
rect 2562 13567 2878 13568
rect 7562 13632 7878 13633
rect 7562 13568 7568 13632
rect 7632 13568 7648 13632
rect 7712 13568 7728 13632
rect 7792 13568 7808 13632
rect 7872 13568 7878 13632
rect 7562 13567 7878 13568
rect 8477 13562 8543 13565
rect 11973 13562 12039 13565
rect 8477 13560 12039 13562
rect 8477 13504 8482 13560
rect 8538 13504 11978 13560
rect 12034 13504 12039 13560
rect 8477 13502 12039 13504
rect 8477 13499 8543 13502
rect 11973 13499 12039 13502
rect 4521 13426 4587 13429
rect 7925 13426 7991 13429
rect 11329 13426 11395 13429
rect 4521 13424 7850 13426
rect 4521 13368 4526 13424
rect 4582 13368 7850 13424
rect 4521 13366 7850 13368
rect 4521 13363 4587 13366
rect 1117 13290 1183 13293
rect 5165 13290 5231 13293
rect 1117 13288 5231 13290
rect 1117 13232 1122 13288
rect 1178 13232 5170 13288
rect 5226 13232 5231 13288
rect 1117 13230 5231 13232
rect 7790 13290 7850 13366
rect 7925 13424 11395 13426
rect 7925 13368 7930 13424
rect 7986 13368 11334 13424
rect 11390 13368 11395 13424
rect 14000 13392 34000 13512
rect 7925 13366 11395 13368
rect 7925 13363 7991 13366
rect 11329 13363 11395 13366
rect 16622 13293 16682 13392
rect 9121 13290 9187 13293
rect 12709 13290 12775 13293
rect 16297 13290 16363 13293
rect 7790 13230 9000 13290
rect 1117 13227 1183 13230
rect 5165 13227 5231 13230
rect 8940 13154 9000 13230
rect 9121 13288 12775 13290
rect 9121 13232 9126 13288
rect 9182 13232 12714 13288
rect 12770 13232 12775 13288
rect 9121 13230 12775 13232
rect 9121 13227 9187 13230
rect 12709 13227 12775 13230
rect 13310 13288 16363 13290
rect 13310 13232 16302 13288
rect 16358 13232 16363 13288
rect 13310 13230 16363 13232
rect 16622 13288 16731 13293
rect 16622 13232 16670 13288
rect 16726 13232 16731 13288
rect 16622 13230 16731 13232
rect 10961 13154 11027 13157
rect 8940 13152 11027 13154
rect 8940 13096 10966 13152
rect 11022 13096 11027 13152
rect 8940 13094 11027 13096
rect 10961 13091 11027 13094
rect 3562 13088 3878 13089
rect 3562 13024 3568 13088
rect 3632 13024 3648 13088
rect 3712 13024 3728 13088
rect 3792 13024 3808 13088
rect 3872 13024 3878 13088
rect 3562 13023 3878 13024
rect 8562 13088 8878 13089
rect 8562 13024 8568 13088
rect 8632 13024 8648 13088
rect 8712 13024 8728 13088
rect 8792 13024 8808 13088
rect 8872 13024 8878 13088
rect 8562 13023 8878 13024
rect 1577 13018 1643 13021
rect 3049 13018 3115 13021
rect 1577 13016 3115 13018
rect 1577 12960 1582 13016
rect 1638 12960 3054 13016
rect 3110 12960 3115 13016
rect 1577 12958 3115 12960
rect 1577 12955 1643 12958
rect 3049 12955 3115 12958
rect 9029 13018 9095 13021
rect 13310 13018 13370 13230
rect 16297 13227 16363 13230
rect 16665 13227 16731 13230
rect 9029 13016 13370 13018
rect 9029 12960 9034 13016
rect 9090 12960 13370 13016
rect 9029 12958 13370 12960
rect 13445 13018 13511 13021
rect 14000 13018 34000 13104
rect 13445 13016 34000 13018
rect 13445 12960 13450 13016
rect 13506 12984 34000 13016
rect 13506 12960 14076 12984
rect 13445 12958 14076 12960
rect 9029 12955 9095 12958
rect 13445 12955 13511 12958
rect 1485 12882 1551 12885
rect 3417 12882 3483 12885
rect 1485 12880 3483 12882
rect 1485 12824 1490 12880
rect 1546 12824 3422 12880
rect 3478 12824 3483 12880
rect 1485 12822 3483 12824
rect 1485 12819 1551 12822
rect 3417 12819 3483 12822
rect 3877 12882 3943 12885
rect 8017 12882 8083 12885
rect 3877 12880 8083 12882
rect 3877 12824 3882 12880
rect 3938 12824 8022 12880
rect 8078 12824 8083 12880
rect 3877 12822 8083 12824
rect 3877 12819 3943 12822
rect 8017 12819 8083 12822
rect 8201 12882 8267 12885
rect 12525 12882 12591 12885
rect 8201 12880 12591 12882
rect 8201 12824 8206 12880
rect 8262 12824 12530 12880
rect 12586 12824 12591 12880
rect 8201 12822 12591 12824
rect 8201 12819 8267 12822
rect 12525 12819 12591 12822
rect 2262 12684 2268 12748
rect 2332 12746 2338 12748
rect 2497 12746 2563 12749
rect 2332 12744 2563 12746
rect 2332 12688 2502 12744
rect 2558 12688 2563 12744
rect 2332 12686 2563 12688
rect 2332 12684 2338 12686
rect 2497 12683 2563 12686
rect 6637 12746 6703 12749
rect 13813 12746 13879 12749
rect 6637 12744 13879 12746
rect 6637 12688 6642 12744
rect 6698 12688 13818 12744
rect 13874 12688 13879 12744
rect 6637 12686 13879 12688
rect 6637 12683 6703 12686
rect 13813 12683 13879 12686
rect 7281 12610 7347 12613
rect 4064 12608 7347 12610
rect 4064 12552 7286 12608
rect 7342 12552 7347 12608
rect 4064 12550 7347 12552
rect 2562 12544 2878 12545
rect 2562 12480 2568 12544
rect 2632 12480 2648 12544
rect 2712 12480 2728 12544
rect 2792 12480 2808 12544
rect 2872 12480 2878 12544
rect 2562 12479 2878 12480
rect 4064 12477 4124 12550
rect 7281 12547 7347 12550
rect 8017 12610 8083 12613
rect 13721 12610 13787 12613
rect 8017 12608 13787 12610
rect 8017 12552 8022 12608
rect 8078 12552 13726 12608
rect 13782 12552 13787 12608
rect 14000 12576 34000 12696
rect 8017 12550 13787 12552
rect 8017 12547 8083 12550
rect 13721 12547 13787 12550
rect 7562 12544 7878 12545
rect 7562 12480 7568 12544
rect 7632 12480 7648 12544
rect 7712 12480 7728 12544
rect 7792 12480 7808 12544
rect 7872 12480 7878 12544
rect 7562 12479 7878 12480
rect 15886 12477 15946 12576
rect 3233 12474 3299 12477
rect 4061 12474 4127 12477
rect 3233 12472 4127 12474
rect 3233 12416 3238 12472
rect 3294 12416 4066 12472
rect 4122 12416 4127 12472
rect 3233 12414 4127 12416
rect 3233 12411 3299 12414
rect 4061 12411 4127 12414
rect 4337 12474 4403 12477
rect 8937 12474 9003 12477
rect 4337 12472 7482 12474
rect 4337 12416 4342 12472
rect 4398 12416 7482 12472
rect 4337 12414 7482 12416
rect 4337 12411 4403 12414
rect 2681 12338 2747 12341
rect 4061 12338 4127 12341
rect 5717 12338 5783 12341
rect 2681 12336 4127 12338
rect 2681 12280 2686 12336
rect 2742 12280 4066 12336
rect 4122 12280 4127 12336
rect 2681 12278 4127 12280
rect 2681 12275 2747 12278
rect 4061 12275 4127 12278
rect 4478 12336 5783 12338
rect 4478 12280 5722 12336
rect 5778 12280 5783 12336
rect 4478 12278 5783 12280
rect 7422 12338 7482 12414
rect 7974 12472 9003 12474
rect 7974 12416 8942 12472
rect 8998 12416 9003 12472
rect 7974 12414 9003 12416
rect 7974 12338 8034 12414
rect 8937 12411 9003 12414
rect 9213 12474 9279 12477
rect 15653 12474 15719 12477
rect 9213 12472 15719 12474
rect 9213 12416 9218 12472
rect 9274 12416 15658 12472
rect 15714 12416 15719 12472
rect 9213 12414 15719 12416
rect 15886 12472 15995 12477
rect 15886 12416 15934 12472
rect 15990 12416 15995 12472
rect 15886 12414 15995 12416
rect 9213 12411 9279 12414
rect 7422 12278 8034 12338
rect 2313 12202 2379 12205
rect 4337 12202 4403 12205
rect 2313 12200 4403 12202
rect 2313 12144 2318 12200
rect 2374 12144 4342 12200
rect 4398 12144 4403 12200
rect 2313 12142 4403 12144
rect 2313 12139 2379 12142
rect 4337 12139 4403 12142
rect 3969 12066 4035 12069
rect 4478 12066 4538 12278
rect 5717 12275 5783 12278
rect 4981 12202 5047 12205
rect 5993 12202 6059 12205
rect 8937 12202 9003 12205
rect 4981 12200 9003 12202
rect 4981 12144 4986 12200
rect 5042 12144 5998 12200
rect 6054 12144 8942 12200
rect 8998 12144 9003 12200
rect 4981 12142 9003 12144
rect 4981 12139 5047 12142
rect 5993 12139 6059 12142
rect 8937 12139 9003 12142
rect 11605 12202 11671 12205
rect 13261 12202 13327 12205
rect 11605 12200 13327 12202
rect 11605 12144 11610 12200
rect 11666 12144 13266 12200
rect 13322 12144 13327 12200
rect 11605 12142 13327 12144
rect 13862 12202 13922 12414
rect 15653 12411 15719 12414
rect 15929 12411 15995 12414
rect 14000 12202 34000 12288
rect 13862 12168 34000 12202
rect 13862 12142 14076 12168
rect 11605 12139 11671 12142
rect 13261 12139 13327 12142
rect 3969 12064 4538 12066
rect 3969 12008 3974 12064
rect 4030 12008 4538 12064
rect 3969 12006 4538 12008
rect 3969 12003 4035 12006
rect 9254 12004 9260 12068
rect 9324 12066 9330 12068
rect 15285 12066 15351 12069
rect 9324 12064 15351 12066
rect 9324 12008 15290 12064
rect 15346 12008 15351 12064
rect 9324 12006 15351 12008
rect 9324 12004 9330 12006
rect 15285 12003 15351 12006
rect 3562 12000 3878 12001
rect 3562 11936 3568 12000
rect 3632 11936 3648 12000
rect 3712 11936 3728 12000
rect 3792 11936 3808 12000
rect 3872 11936 3878 12000
rect 3562 11935 3878 11936
rect 8562 12000 8878 12001
rect 8562 11936 8568 12000
rect 8632 11936 8648 12000
rect 8712 11936 8728 12000
rect 8792 11936 8808 12000
rect 8872 11936 8878 12000
rect 8562 11935 8878 11936
rect 6821 11794 6887 11797
rect 11329 11794 11395 11797
rect 6821 11792 11395 11794
rect 6821 11736 6826 11792
rect 6882 11736 11334 11792
rect 11390 11736 11395 11792
rect 14000 11760 34000 11880
rect 6821 11734 11395 11736
rect 6821 11731 6887 11734
rect 11329 11731 11395 11734
rect 15334 11661 15394 11760
rect 7189 11658 7255 11661
rect 13445 11658 13511 11661
rect 7189 11656 13511 11658
rect 7189 11600 7194 11656
rect 7250 11600 13450 11656
rect 13506 11600 13511 11656
rect 7189 11598 13511 11600
rect 15334 11656 15443 11661
rect 15334 11600 15382 11656
rect 15438 11600 15443 11656
rect 15334 11598 15443 11600
rect 7189 11595 7255 11598
rect 13445 11595 13511 11598
rect 15377 11595 15443 11598
rect 11973 11522 12039 11525
rect 12617 11522 12683 11525
rect 11973 11520 12683 11522
rect 11973 11464 11978 11520
rect 12034 11464 12622 11520
rect 12678 11464 12683 11520
rect 11973 11462 12683 11464
rect 11973 11459 12039 11462
rect 12617 11459 12683 11462
rect 2562 11456 2878 11457
rect 2562 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2878 11456
rect 2562 11391 2878 11392
rect 7562 11456 7878 11457
rect 7562 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7878 11456
rect 7562 11391 7878 11392
rect 9029 11386 9095 11389
rect 8020 11384 9095 11386
rect 8020 11328 9034 11384
rect 9090 11328 9095 11384
rect 8020 11326 9095 11328
rect 4153 11250 4219 11253
rect 8020 11250 8080 11326
rect 9029 11323 9095 11326
rect 9213 11386 9279 11389
rect 12341 11386 12407 11389
rect 9213 11384 12407 11386
rect 9213 11328 9218 11384
rect 9274 11328 12346 11384
rect 12402 11328 12407 11384
rect 9213 11326 12407 11328
rect 9213 11323 9279 11326
rect 12341 11323 12407 11326
rect 12525 11386 12591 11389
rect 14000 11386 34000 11472
rect 12525 11384 34000 11386
rect 12525 11328 12530 11384
rect 12586 11352 34000 11384
rect 12586 11328 14076 11352
rect 12525 11326 14076 11328
rect 12525 11323 12591 11326
rect 4153 11248 8080 11250
rect 4153 11192 4158 11248
rect 4214 11192 8080 11248
rect 4153 11190 8080 11192
rect 8201 11250 8267 11253
rect 11145 11250 11211 11253
rect 8201 11248 11211 11250
rect 8201 11192 8206 11248
rect 8262 11192 11150 11248
rect 11206 11192 11211 11248
rect 8201 11190 11211 11192
rect 4153 11187 4219 11190
rect 8201 11187 8267 11190
rect 11145 11187 11211 11190
rect 11329 11250 11395 11253
rect 12893 11250 12959 11253
rect 15377 11250 15443 11253
rect 11329 11248 12959 11250
rect 11329 11192 11334 11248
rect 11390 11192 12898 11248
rect 12954 11192 12959 11248
rect 11329 11190 12959 11192
rect 11329 11187 11395 11190
rect 12893 11187 12959 11190
rect 13862 11248 15443 11250
rect 13862 11192 15382 11248
rect 15438 11192 15443 11248
rect 13862 11190 15443 11192
rect 5165 11114 5231 11117
rect 7097 11114 7163 11117
rect 5165 11112 7163 11114
rect 5165 11056 5170 11112
rect 5226 11056 7102 11112
rect 7158 11056 7163 11112
rect 5165 11054 7163 11056
rect 5165 11051 5231 11054
rect 7097 11051 7163 11054
rect 9121 11114 9187 11117
rect 13862 11114 13922 11190
rect 15377 11187 15443 11190
rect 9121 11112 13922 11114
rect 9121 11056 9126 11112
rect 9182 11056 13922 11112
rect 9121 11054 13922 11056
rect 9121 11051 9187 11054
rect 14000 10944 34000 11064
rect 3562 10912 3878 10913
rect 3562 10848 3568 10912
rect 3632 10848 3648 10912
rect 3712 10848 3728 10912
rect 3792 10848 3808 10912
rect 3872 10848 3878 10912
rect 3562 10847 3878 10848
rect 8562 10912 8878 10913
rect 8562 10848 8568 10912
rect 8632 10848 8648 10912
rect 8712 10848 8728 10912
rect 8792 10848 8808 10912
rect 8872 10848 8878 10912
rect 8562 10847 8878 10848
rect 16438 10845 16498 10944
rect 13629 10842 13695 10845
rect 16113 10842 16179 10845
rect 13629 10840 16179 10842
rect 13629 10784 13634 10840
rect 13690 10784 16118 10840
rect 16174 10784 16179 10840
rect 13629 10782 16179 10784
rect 13629 10779 13695 10782
rect 16113 10779 16179 10782
rect 16389 10840 16498 10845
rect 16389 10784 16394 10840
rect 16450 10784 16498 10840
rect 16389 10782 16498 10784
rect 16389 10779 16455 10782
rect 197 10706 263 10709
rect 2221 10706 2287 10709
rect 197 10704 2287 10706
rect 197 10648 202 10704
rect 258 10648 2226 10704
rect 2282 10648 2287 10704
rect 197 10646 2287 10648
rect 197 10643 263 10646
rect 2221 10643 2287 10646
rect 2405 10706 2471 10709
rect 5257 10706 5323 10709
rect 5625 10706 5691 10709
rect 2405 10704 5691 10706
rect 2405 10648 2410 10704
rect 2466 10648 5262 10704
rect 5318 10648 5630 10704
rect 5686 10648 5691 10704
rect 2405 10646 5691 10648
rect 2405 10643 2471 10646
rect 5257 10643 5323 10646
rect 5625 10643 5691 10646
rect 11053 10706 11119 10709
rect 12525 10706 12591 10709
rect 11053 10704 12591 10706
rect 11053 10648 11058 10704
rect 11114 10648 12530 10704
rect 12586 10648 12591 10704
rect 11053 10646 12591 10648
rect 11053 10643 11119 10646
rect 12525 10643 12591 10646
rect 12709 10706 12775 10709
rect 12709 10704 13692 10706
rect 12709 10648 12714 10704
rect 12770 10648 13692 10704
rect 12709 10646 13692 10648
rect 12709 10643 12775 10646
rect 5349 10570 5415 10573
rect 13445 10570 13511 10573
rect 5349 10568 13511 10570
rect 5349 10512 5354 10568
rect 5410 10512 13450 10568
rect 13506 10512 13511 10568
rect 5349 10510 13511 10512
rect 13632 10570 13692 10646
rect 14000 10570 34000 10656
rect 13632 10536 34000 10570
rect 13632 10510 14076 10536
rect 5349 10507 5415 10510
rect 13445 10507 13511 10510
rect 9213 10434 9279 10437
rect 13905 10434 13971 10437
rect 9213 10432 13971 10434
rect 9213 10376 9218 10432
rect 9274 10376 13910 10432
rect 13966 10376 13971 10432
rect 9213 10374 13971 10376
rect 9213 10371 9279 10374
rect 13905 10371 13971 10374
rect 14365 10434 14431 10437
rect 15561 10434 15627 10437
rect 14365 10432 15627 10434
rect 14365 10376 14370 10432
rect 14426 10376 15566 10432
rect 15622 10376 15627 10432
rect 14365 10374 15627 10376
rect 14365 10371 14431 10374
rect 15561 10371 15627 10374
rect 2562 10368 2878 10369
rect 2562 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2878 10368
rect 2562 10303 2878 10304
rect 7562 10368 7878 10369
rect 7562 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7878 10368
rect 7562 10303 7878 10304
rect 4061 10162 4127 10165
rect 5993 10162 6059 10165
rect 4061 10160 6059 10162
rect 4061 10104 4066 10160
rect 4122 10104 5998 10160
rect 6054 10104 6059 10160
rect 4061 10102 6059 10104
rect 4061 10099 4127 10102
rect 5993 10099 6059 10102
rect 13813 10162 13879 10165
rect 14000 10162 34000 10248
rect 13813 10160 34000 10162
rect 13813 10104 13818 10160
rect 13874 10128 34000 10160
rect 13874 10104 14076 10128
rect 13813 10102 14076 10104
rect 13813 10099 13879 10102
rect 8017 10026 8083 10029
rect 12709 10026 12775 10029
rect 8017 10024 12775 10026
rect 8017 9968 8022 10024
rect 8078 9968 12714 10024
rect 12770 9968 12775 10024
rect 8017 9966 12775 9968
rect 8017 9963 8083 9966
rect 12709 9963 12775 9966
rect 9857 9890 9923 9893
rect 13077 9890 13143 9893
rect 9857 9888 13143 9890
rect 9857 9832 9862 9888
rect 9918 9832 13082 9888
rect 13138 9832 13143 9888
rect 9857 9830 13143 9832
rect 9857 9827 9923 9830
rect 13077 9827 13143 9830
rect 3562 9824 3878 9825
rect 3562 9760 3568 9824
rect 3632 9760 3648 9824
rect 3712 9760 3728 9824
rect 3792 9760 3808 9824
rect 3872 9760 3878 9824
rect 3562 9759 3878 9760
rect 8562 9824 8878 9825
rect 8562 9760 8568 9824
rect 8632 9760 8648 9824
rect 8712 9760 8728 9824
rect 8792 9760 8808 9824
rect 8872 9760 8878 9824
rect 8562 9759 8878 9760
rect 5349 9754 5415 9757
rect 8385 9754 8451 9757
rect 5349 9752 8451 9754
rect 5349 9696 5354 9752
rect 5410 9696 8390 9752
rect 8446 9696 8451 9752
rect 5349 9694 8451 9696
rect 5349 9691 5415 9694
rect 8385 9691 8451 9694
rect 11145 9754 11211 9757
rect 12801 9754 12867 9757
rect 11145 9752 12867 9754
rect 11145 9696 11150 9752
rect 11206 9696 12806 9752
rect 12862 9696 12867 9752
rect 11145 9694 12867 9696
rect 11145 9691 11211 9694
rect 12801 9691 12867 9694
rect 13721 9754 13787 9757
rect 14000 9754 34000 9840
rect 13721 9752 34000 9754
rect 13721 9696 13726 9752
rect 13782 9720 34000 9752
rect 13782 9696 14076 9720
rect 13721 9694 14076 9696
rect 13721 9691 13787 9694
rect 1945 9618 2011 9621
rect 5441 9618 5507 9621
rect 1945 9616 5507 9618
rect 1945 9560 1950 9616
rect 2006 9560 5446 9616
rect 5502 9560 5507 9616
rect 1945 9558 5507 9560
rect 1945 9555 2011 9558
rect 5441 9555 5507 9558
rect 5809 9618 5875 9621
rect 8477 9618 8543 9621
rect 5809 9616 8543 9618
rect 5809 9560 5814 9616
rect 5870 9560 8482 9616
rect 8538 9560 8543 9616
rect 5809 9558 8543 9560
rect 5809 9555 5875 9558
rect 8477 9555 8543 9558
rect 9121 9618 9187 9621
rect 15193 9618 15259 9621
rect 9121 9616 15259 9618
rect 9121 9560 9126 9616
rect 9182 9560 15198 9616
rect 15254 9560 15259 9616
rect 9121 9558 15259 9560
rect 9121 9555 9187 9558
rect 15193 9555 15259 9558
rect 6821 9482 6887 9485
rect 9305 9482 9371 9485
rect 6821 9480 9371 9482
rect 6821 9424 6826 9480
rect 6882 9424 9310 9480
rect 9366 9424 9371 9480
rect 6821 9422 9371 9424
rect 6821 9419 6887 9422
rect 9305 9419 9371 9422
rect 13813 9346 13879 9349
rect 14000 9346 34000 9432
rect 13813 9344 34000 9346
rect 13813 9288 13818 9344
rect 13874 9312 34000 9344
rect 13874 9288 14076 9312
rect 13813 9286 14076 9288
rect 13813 9283 13879 9286
rect 2562 9280 2878 9281
rect 2562 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2878 9280
rect 2562 9215 2878 9216
rect 7562 9280 7878 9281
rect 7562 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7878 9280
rect 7562 9215 7878 9216
rect 8201 9210 8267 9213
rect 13813 9210 13879 9213
rect 8201 9208 13879 9210
rect 8201 9152 8206 9208
rect 8262 9152 13818 9208
rect 13874 9152 13879 9208
rect 8201 9150 13879 9152
rect 8201 9147 8267 9150
rect 13813 9147 13879 9150
rect 4153 9074 4219 9077
rect 5993 9074 6059 9077
rect 4153 9072 6059 9074
rect 4153 9016 4158 9072
rect 4214 9016 5998 9072
rect 6054 9016 6059 9072
rect 4153 9014 6059 9016
rect 4153 9011 4219 9014
rect 5993 9011 6059 9014
rect 6729 9074 6795 9077
rect 9949 9074 10015 9077
rect 6729 9072 10015 9074
rect 6729 9016 6734 9072
rect 6790 9016 9954 9072
rect 10010 9016 10015 9072
rect 6729 9014 10015 9016
rect 6729 9011 6795 9014
rect 9949 9011 10015 9014
rect 5625 8938 5691 8941
rect 11421 8938 11487 8941
rect 5625 8936 11487 8938
rect 5625 8880 5630 8936
rect 5686 8880 11426 8936
rect 11482 8880 11487 8936
rect 5625 8878 11487 8880
rect 5625 8875 5691 8878
rect 11421 8875 11487 8878
rect 13537 8938 13603 8941
rect 14000 8938 34000 9024
rect 13537 8936 34000 8938
rect 13537 8880 13542 8936
rect 13598 8904 34000 8936
rect 13598 8880 14076 8904
rect 13537 8878 14076 8880
rect 13537 8875 13603 8878
rect 9581 8802 9647 8805
rect 13721 8802 13787 8805
rect 9581 8800 13787 8802
rect 9581 8744 9586 8800
rect 9642 8744 13726 8800
rect 13782 8744 13787 8800
rect 9581 8742 13787 8744
rect 9581 8739 9647 8742
rect 13721 8739 13787 8742
rect 3562 8736 3878 8737
rect 3562 8672 3568 8736
rect 3632 8672 3648 8736
rect 3712 8672 3728 8736
rect 3792 8672 3808 8736
rect 3872 8672 3878 8736
rect 3562 8671 3878 8672
rect 8562 8736 8878 8737
rect 8562 8672 8568 8736
rect 8632 8672 8648 8736
rect 8712 8672 8728 8736
rect 8792 8672 8808 8736
rect 8872 8672 8878 8736
rect 8562 8671 8878 8672
rect 3969 8666 4035 8669
rect 5257 8666 5323 8669
rect 3969 8664 5323 8666
rect 3969 8608 3974 8664
rect 4030 8608 5262 8664
rect 5318 8608 5323 8664
rect 3969 8606 5323 8608
rect 3969 8603 4035 8606
rect 5257 8603 5323 8606
rect 3141 8530 3207 8533
rect 6361 8530 6427 8533
rect 3141 8528 6427 8530
rect 3141 8472 3146 8528
rect 3202 8472 6366 8528
rect 6422 8472 6427 8528
rect 3141 8470 6427 8472
rect 3141 8467 3207 8470
rect 6361 8467 6427 8470
rect 6821 8530 6887 8533
rect 14000 8530 34000 8616
rect 6821 8528 34000 8530
rect 6821 8472 6826 8528
rect 6882 8496 34000 8528
rect 6882 8472 14076 8496
rect 6821 8470 14076 8472
rect 6821 8467 6887 8470
rect 1761 8394 1827 8397
rect 3417 8394 3483 8397
rect 1761 8392 3483 8394
rect 1761 8336 1766 8392
rect 1822 8336 3422 8392
rect 3478 8336 3483 8392
rect 1761 8334 3483 8336
rect 1761 8331 1827 8334
rect 3417 8331 3483 8334
rect 13077 8394 13143 8397
rect 13997 8394 14063 8397
rect 13077 8392 14063 8394
rect 13077 8336 13082 8392
rect 13138 8336 14002 8392
rect 14058 8336 14063 8392
rect 13077 8334 14063 8336
rect 13077 8331 13143 8334
rect 13997 8331 14063 8334
rect 15561 8394 15627 8397
rect 16481 8394 16547 8397
rect 15561 8392 16547 8394
rect 15561 8336 15566 8392
rect 15622 8336 16486 8392
rect 16542 8336 16547 8392
rect 15561 8334 16547 8336
rect 15561 8331 15627 8334
rect 16481 8331 16547 8334
rect 6862 8196 6868 8260
rect 6932 8258 6938 8260
rect 7189 8258 7255 8261
rect 6932 8256 7255 8258
rect 6932 8200 7194 8256
rect 7250 8200 7255 8256
rect 6932 8198 7255 8200
rect 6932 8196 6938 8198
rect 7189 8195 7255 8198
rect 9857 8258 9923 8261
rect 12525 8258 12591 8261
rect 9857 8256 12591 8258
rect 9857 8200 9862 8256
rect 9918 8200 12530 8256
rect 12586 8200 12591 8256
rect 9857 8198 12591 8200
rect 9857 8195 9923 8198
rect 12525 8195 12591 8198
rect 2562 8192 2878 8193
rect 2562 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2878 8192
rect 2562 8127 2878 8128
rect 7562 8192 7878 8193
rect 7562 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7878 8192
rect 7562 8127 7878 8128
rect 13721 8122 13787 8125
rect 14000 8122 34000 8208
rect 13721 8120 34000 8122
rect 13721 8064 13726 8120
rect 13782 8088 34000 8120
rect 13782 8064 14076 8088
rect 13721 8062 14076 8064
rect 13721 8059 13787 8062
rect 2262 7924 2268 7988
rect 2332 7986 2338 7988
rect 15469 7986 15535 7989
rect 2332 7984 15535 7986
rect 2332 7928 15474 7984
rect 15530 7928 15535 7984
rect 2332 7926 15535 7928
rect 2332 7924 2338 7926
rect 15469 7923 15535 7926
rect 2129 7850 2195 7853
rect 2129 7848 5826 7850
rect 2129 7792 2134 7848
rect 2190 7792 5826 7848
rect 2129 7790 5826 7792
rect 2129 7787 2195 7790
rect 5766 7714 5826 7790
rect 8293 7714 8359 7717
rect 5766 7712 8359 7714
rect 5766 7656 8298 7712
rect 8354 7656 8359 7712
rect 5766 7654 8359 7656
rect 8293 7651 8359 7654
rect 11789 7714 11855 7717
rect 14000 7714 34000 7800
rect 11789 7712 34000 7714
rect 11789 7656 11794 7712
rect 11850 7680 34000 7712
rect 11850 7656 14076 7680
rect 11789 7654 14076 7656
rect 11789 7651 11855 7654
rect 3562 7648 3878 7649
rect 3562 7584 3568 7648
rect 3632 7584 3648 7648
rect 3712 7584 3728 7648
rect 3792 7584 3808 7648
rect 3872 7584 3878 7648
rect 3562 7583 3878 7584
rect 8562 7648 8878 7649
rect 8562 7584 8568 7648
rect 8632 7584 8648 7648
rect 8712 7584 8728 7648
rect 8792 7584 8808 7648
rect 8872 7584 8878 7648
rect 8562 7583 8878 7584
rect 5901 7578 5967 7581
rect 7097 7578 7163 7581
rect 5901 7576 7163 7578
rect 5901 7520 5906 7576
rect 5962 7520 7102 7576
rect 7158 7520 7163 7576
rect 5901 7518 7163 7520
rect 5901 7515 5967 7518
rect 7097 7515 7163 7518
rect 13905 7578 13971 7581
rect 15929 7578 15995 7581
rect 13905 7576 15995 7578
rect 13905 7520 13910 7576
rect 13966 7520 15934 7576
rect 15990 7520 15995 7576
rect 13905 7518 15995 7520
rect 13905 7515 13971 7518
rect 15929 7515 15995 7518
rect 4981 7306 5047 7309
rect 7373 7306 7439 7309
rect 4981 7304 7439 7306
rect 4981 7248 4986 7304
rect 5042 7248 7378 7304
rect 7434 7248 7439 7304
rect 4981 7246 7439 7248
rect 4981 7243 5047 7246
rect 7373 7243 7439 7246
rect 13353 7306 13419 7309
rect 14000 7306 34000 7392
rect 13353 7304 34000 7306
rect 13353 7248 13358 7304
rect 13414 7272 34000 7304
rect 13414 7248 14076 7272
rect 13353 7246 14076 7248
rect 13353 7243 13419 7246
rect 4889 7170 4955 7173
rect 7097 7170 7163 7173
rect 4889 7168 7163 7170
rect 4889 7112 4894 7168
rect 4950 7112 7102 7168
rect 7158 7112 7163 7168
rect 4889 7110 7163 7112
rect 4889 7107 4955 7110
rect 7097 7107 7163 7110
rect 2562 7104 2878 7105
rect 2562 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2878 7104
rect 2562 7039 2878 7040
rect 7562 7104 7878 7105
rect 7562 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7878 7104
rect 7562 7039 7878 7040
rect 2957 7034 3023 7037
rect 6361 7034 6427 7037
rect 2957 7032 6427 7034
rect 2957 6976 2962 7032
rect 3018 6976 6366 7032
rect 6422 6976 6427 7032
rect 2957 6974 6427 6976
rect 2957 6971 3023 6974
rect 6361 6971 6427 6974
rect 6637 6898 6703 6901
rect 13445 6898 13511 6901
rect 6637 6896 13511 6898
rect 6637 6840 6642 6896
rect 6698 6840 13450 6896
rect 13506 6840 13511 6896
rect 6637 6838 13511 6840
rect 6637 6835 6703 6838
rect 13445 6835 13511 6838
rect 13629 6898 13695 6901
rect 14000 6898 34000 6984
rect 13629 6896 34000 6898
rect 13629 6840 13634 6896
rect 13690 6864 34000 6896
rect 13690 6840 14076 6864
rect 13629 6838 14076 6840
rect 13629 6835 13695 6838
rect 5809 6762 5875 6765
rect 13721 6762 13787 6765
rect 15377 6762 15443 6765
rect 5809 6760 13787 6762
rect 5809 6704 5814 6760
rect 5870 6704 13726 6760
rect 13782 6704 13787 6760
rect 5809 6702 13787 6704
rect 5809 6699 5875 6702
rect 13721 6699 13787 6702
rect 13862 6760 15443 6762
rect 13862 6704 15382 6760
rect 15438 6704 15443 6760
rect 13862 6702 15443 6704
rect 12617 6626 12683 6629
rect 8940 6624 12683 6626
rect 8940 6568 12622 6624
rect 12678 6568 12683 6624
rect 8940 6566 12683 6568
rect 3562 6560 3878 6561
rect 3562 6496 3568 6560
rect 3632 6496 3648 6560
rect 3712 6496 3728 6560
rect 3792 6496 3808 6560
rect 3872 6496 3878 6560
rect 3562 6495 3878 6496
rect 8562 6560 8878 6561
rect 8562 6496 8568 6560
rect 8632 6496 8648 6560
rect 8712 6496 8728 6560
rect 8792 6496 8808 6560
rect 8872 6496 8878 6560
rect 8562 6495 8878 6496
rect 2221 6492 2287 6493
rect 2221 6490 2268 6492
rect 2176 6488 2268 6490
rect 2176 6432 2226 6488
rect 2176 6430 2268 6432
rect 2221 6428 2268 6430
rect 2332 6428 2338 6492
rect 2221 6427 2287 6428
rect 8940 6357 9000 6566
rect 12617 6563 12683 6566
rect 13445 6626 13511 6629
rect 13862 6626 13922 6702
rect 15377 6699 15443 6702
rect 13445 6624 13922 6626
rect 13445 6568 13450 6624
rect 13506 6568 13922 6624
rect 13445 6566 13922 6568
rect 13445 6563 13511 6566
rect 10133 6490 10199 6493
rect 14000 6490 34000 6576
rect 10133 6488 34000 6490
rect 10133 6432 10138 6488
rect 10194 6456 34000 6488
rect 10194 6432 14076 6456
rect 10133 6430 14076 6432
rect 10133 6427 10199 6430
rect 5809 6354 5875 6357
rect 8937 6354 9003 6357
rect 5809 6352 9003 6354
rect 5809 6296 5814 6352
rect 5870 6296 8942 6352
rect 8998 6296 9003 6352
rect 5809 6294 9003 6296
rect 5809 6291 5875 6294
rect 8937 6291 9003 6294
rect 9121 6354 9187 6357
rect 13537 6354 13603 6357
rect 9121 6352 13603 6354
rect 9121 6296 9126 6352
rect 9182 6296 13542 6352
rect 13598 6296 13603 6352
rect 9121 6294 13603 6296
rect 9121 6291 9187 6294
rect 13537 6291 13603 6294
rect 13721 6354 13787 6357
rect 16389 6354 16455 6357
rect 13721 6352 16455 6354
rect 13721 6296 13726 6352
rect 13782 6296 16394 6352
rect 16450 6296 16455 6352
rect 13721 6294 16455 6296
rect 13721 6291 13787 6294
rect 16389 6291 16455 6294
rect 1485 6218 1551 6221
rect 13813 6218 13879 6221
rect 1485 6216 13879 6218
rect 1485 6160 1490 6216
rect 1546 6160 13818 6216
rect 13874 6160 13879 6216
rect 1485 6158 13879 6160
rect 1485 6155 1551 6158
rect 13813 6155 13879 6158
rect 5901 6082 5967 6085
rect 3006 6080 5967 6082
rect 3006 6024 5906 6080
rect 5962 6024 5967 6080
rect 3006 6022 5967 6024
rect 2562 6016 2878 6017
rect 2562 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2878 6016
rect 2562 5951 2878 5952
rect 2221 5810 2287 5813
rect 3006 5810 3066 6022
rect 5901 6019 5967 6022
rect 12525 6082 12591 6085
rect 13721 6082 13787 6085
rect 12525 6080 13787 6082
rect 12525 6024 12530 6080
rect 12586 6024 13726 6080
rect 13782 6024 13787 6080
rect 14000 6048 34000 6168
rect 12525 6022 13787 6024
rect 12525 6019 12591 6022
rect 13721 6019 13787 6022
rect 7562 6016 7878 6017
rect 7562 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7878 6016
rect 7562 5951 7878 5952
rect 16622 5949 16682 6048
rect 3233 5946 3299 5949
rect 4521 5946 4587 5949
rect 3233 5944 4587 5946
rect 3233 5888 3238 5944
rect 3294 5888 4526 5944
rect 4582 5888 4587 5944
rect 3233 5886 4587 5888
rect 3233 5883 3299 5886
rect 4521 5883 4587 5886
rect 5073 5946 5139 5949
rect 5717 5946 5783 5949
rect 5073 5944 5783 5946
rect 5073 5888 5078 5944
rect 5134 5888 5722 5944
rect 5778 5888 5783 5944
rect 5073 5886 5783 5888
rect 5073 5883 5139 5886
rect 5717 5883 5783 5886
rect 8201 5946 8267 5949
rect 16481 5946 16547 5949
rect 8201 5944 16547 5946
rect 8201 5888 8206 5944
rect 8262 5888 16486 5944
rect 16542 5888 16547 5944
rect 8201 5886 16547 5888
rect 16622 5944 16731 5949
rect 16622 5888 16670 5944
rect 16726 5888 16731 5944
rect 16622 5886 16731 5888
rect 8201 5883 8267 5886
rect 16481 5883 16547 5886
rect 16665 5883 16731 5886
rect 6821 5810 6887 5813
rect 2221 5808 3066 5810
rect 2221 5752 2226 5808
rect 2282 5752 3066 5808
rect 2221 5750 3066 5752
rect 3190 5808 6887 5810
rect 3190 5752 6826 5808
rect 6882 5752 6887 5808
rect 3190 5750 6887 5752
rect 2221 5747 2287 5750
rect 2589 5674 2655 5677
rect 2589 5672 2882 5674
rect 2589 5616 2594 5672
rect 2650 5616 2882 5672
rect 2589 5614 2882 5616
rect 2589 5611 2655 5614
rect 2822 5538 2882 5614
rect 3190 5538 3250 5750
rect 6821 5747 6887 5750
rect 7281 5810 7347 5813
rect 9857 5810 9923 5813
rect 7281 5808 9923 5810
rect 7281 5752 7286 5808
rect 7342 5752 9862 5808
rect 9918 5752 9923 5808
rect 7281 5750 9923 5752
rect 7281 5747 7347 5750
rect 9857 5747 9923 5750
rect 3509 5674 3575 5677
rect 6269 5674 6335 5677
rect 3509 5672 6335 5674
rect 3509 5616 3514 5672
rect 3570 5616 6274 5672
rect 6330 5616 6335 5672
rect 3509 5614 6335 5616
rect 3509 5611 3575 5614
rect 6269 5611 6335 5614
rect 8201 5674 8267 5677
rect 9489 5674 9555 5677
rect 8201 5672 9555 5674
rect 8201 5616 8206 5672
rect 8262 5616 9494 5672
rect 9550 5616 9555 5672
rect 8201 5614 9555 5616
rect 8201 5611 8267 5614
rect 9489 5611 9555 5614
rect 13813 5674 13879 5677
rect 14000 5674 34000 5760
rect 13813 5672 34000 5674
rect 13813 5616 13818 5672
rect 13874 5640 34000 5672
rect 13874 5616 14076 5640
rect 13813 5614 14076 5616
rect 13813 5611 13879 5614
rect 2822 5478 3250 5538
rect 4061 5538 4127 5541
rect 6862 5538 6868 5540
rect 4061 5536 6868 5538
rect 4061 5480 4066 5536
rect 4122 5480 6868 5536
rect 4061 5478 6868 5480
rect 4061 5475 4127 5478
rect 6862 5476 6868 5478
rect 6932 5476 6938 5540
rect 13770 5538 14060 5550
rect 15561 5538 15627 5541
rect 12390 5536 15627 5538
rect 12390 5490 15566 5536
rect 12390 5478 13830 5490
rect 14000 5480 15566 5490
rect 15622 5480 15627 5536
rect 14000 5478 15627 5480
rect 3562 5472 3878 5473
rect 3562 5408 3568 5472
rect 3632 5408 3648 5472
rect 3712 5408 3728 5472
rect 3792 5408 3808 5472
rect 3872 5408 3878 5472
rect 3562 5407 3878 5408
rect 8562 5472 8878 5473
rect 8562 5408 8568 5472
rect 8632 5408 8648 5472
rect 8712 5408 8728 5472
rect 8792 5408 8808 5472
rect 8872 5408 8878 5472
rect 8562 5407 8878 5408
rect 4797 5402 4863 5405
rect 6545 5402 6611 5405
rect 4797 5400 6611 5402
rect 4797 5344 4802 5400
rect 4858 5344 6550 5400
rect 6606 5344 6611 5400
rect 4797 5342 6611 5344
rect 4797 5339 4863 5342
rect 6545 5339 6611 5342
rect 4889 5266 4955 5269
rect 12390 5266 12450 5478
rect 15561 5475 15627 5478
rect 4889 5264 12450 5266
rect 4889 5208 4894 5264
rect 4950 5208 12450 5264
rect 4889 5206 12450 5208
rect 12985 5266 13051 5269
rect 14000 5266 34000 5352
rect 12985 5264 34000 5266
rect 12985 5208 12990 5264
rect 13046 5232 34000 5264
rect 13046 5208 14076 5232
rect 12985 5206 14076 5208
rect 4889 5203 4955 5206
rect 12985 5203 13051 5206
rect 3693 5130 3759 5133
rect 13813 5130 13879 5133
rect 3693 5128 13879 5130
rect 3693 5072 3698 5128
rect 3754 5072 13818 5128
rect 13874 5072 13879 5128
rect 3693 5070 13879 5072
rect 3693 5067 3759 5070
rect 13813 5067 13879 5070
rect 4061 4994 4127 4997
rect 5625 4994 5691 4997
rect 4061 4992 5691 4994
rect 4061 4936 4066 4992
rect 4122 4936 5630 4992
rect 5686 4936 5691 4992
rect 4061 4934 5691 4936
rect 4061 4931 4127 4934
rect 5625 4931 5691 4934
rect 7562 4928 7878 4929
rect 7562 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7878 4928
rect 7562 4863 7878 4864
rect 8385 4858 8451 4861
rect 13629 4858 13695 4861
rect 8385 4856 13695 4858
rect 8385 4800 8390 4856
rect 8446 4800 13634 4856
rect 13690 4800 13695 4856
rect 8385 4798 13695 4800
rect 8385 4795 8451 4798
rect 13629 4795 13695 4798
rect 13813 4858 13879 4861
rect 14000 4858 34000 4944
rect 13813 4856 34000 4858
rect 13813 4800 13818 4856
rect 13874 4824 34000 4856
rect 13874 4800 14076 4824
rect 13813 4798 14076 4800
rect 13813 4795 13879 4798
rect 1669 4722 1735 4725
rect 3325 4722 3391 4725
rect 8569 4722 8635 4725
rect 1669 4720 3391 4722
rect 1669 4664 1674 4720
rect 1730 4664 3330 4720
rect 3386 4664 3391 4720
rect 1669 4662 3391 4664
rect 1669 4659 1735 4662
rect 3325 4659 3391 4662
rect 3558 4720 8635 4722
rect 3558 4664 8574 4720
rect 8630 4664 8635 4720
rect 3558 4662 8635 4664
rect 3141 4586 3207 4589
rect 3558 4586 3618 4662
rect 8569 4659 8635 4662
rect 9305 4722 9371 4725
rect 11421 4722 11487 4725
rect 9305 4720 11487 4722
rect 9305 4664 9310 4720
rect 9366 4664 11426 4720
rect 11482 4664 11487 4720
rect 9305 4662 11487 4664
rect 9305 4659 9371 4662
rect 11421 4659 11487 4662
rect 13905 4722 13971 4725
rect 15101 4722 15167 4725
rect 13905 4720 15167 4722
rect 13905 4664 13910 4720
rect 13966 4664 15106 4720
rect 15162 4664 15167 4720
rect 13905 4662 15167 4664
rect 13905 4659 13971 4662
rect 15101 4659 15167 4662
rect 3141 4584 3618 4586
rect 3141 4528 3146 4584
rect 3202 4528 3618 4584
rect 3141 4526 3618 4528
rect 6913 4586 6979 4589
rect 12341 4586 12407 4589
rect 6913 4584 12407 4586
rect 6913 4528 6918 4584
rect 6974 4528 12346 4584
rect 12402 4528 12407 4584
rect 6913 4526 12407 4528
rect 3141 4523 3207 4526
rect 6913 4523 6979 4526
rect 12341 4523 12407 4526
rect 5625 4450 5691 4453
rect 8385 4450 8451 4453
rect 5625 4448 8451 4450
rect 5625 4392 5630 4448
rect 5686 4392 8390 4448
rect 8446 4392 8451 4448
rect 5625 4390 8451 4392
rect 5625 4387 5691 4390
rect 8385 4387 8451 4390
rect 11881 4450 11947 4453
rect 14000 4450 34000 4536
rect 11881 4448 34000 4450
rect 11881 4392 11886 4448
rect 11942 4416 34000 4448
rect 11942 4392 14076 4416
rect 11881 4390 14076 4392
rect 11881 4387 11947 4390
rect 3562 4384 3878 4385
rect 3562 4320 3568 4384
rect 3632 4320 3648 4384
rect 3712 4320 3728 4384
rect 3792 4320 3808 4384
rect 3872 4320 3878 4384
rect 3562 4319 3878 4320
rect 8562 4384 8878 4385
rect 8562 4320 8568 4384
rect 8632 4320 8648 4384
rect 8712 4320 8728 4384
rect 8792 4320 8808 4384
rect 8872 4320 8878 4384
rect 8562 4319 8878 4320
rect 6085 4314 6151 4317
rect 9305 4314 9371 4317
rect 13997 4314 14063 4317
rect 6085 4312 8218 4314
rect 6085 4256 6090 4312
rect 6146 4256 8218 4312
rect 6085 4254 8218 4256
rect 6085 4251 6151 4254
rect 3049 4178 3115 4181
rect 4337 4178 4403 4181
rect 3049 4176 4403 4178
rect 3049 4120 3054 4176
rect 3110 4120 4342 4176
rect 4398 4120 4403 4176
rect 3049 4118 4403 4120
rect 3049 4115 3115 4118
rect 4337 4115 4403 4118
rect 6269 4178 6335 4181
rect 7925 4178 7991 4181
rect 6269 4176 7991 4178
rect 6269 4120 6274 4176
rect 6330 4120 7930 4176
rect 7986 4120 7991 4176
rect 6269 4118 7991 4120
rect 8158 4178 8218 4254
rect 9305 4312 14063 4314
rect 9305 4256 9310 4312
rect 9366 4256 14002 4312
rect 14058 4256 14063 4312
rect 9305 4254 14063 4256
rect 9305 4251 9371 4254
rect 13997 4251 14063 4254
rect 10961 4178 11027 4181
rect 8158 4176 11027 4178
rect 8158 4120 10966 4176
rect 11022 4120 11027 4176
rect 8158 4118 11027 4120
rect 6269 4115 6335 4118
rect 7925 4115 7991 4118
rect 10961 4115 11027 4118
rect 12433 4178 12499 4181
rect 15837 4178 15903 4181
rect 12433 4176 15903 4178
rect 12433 4120 12438 4176
rect 12494 4120 15842 4176
rect 15898 4120 15903 4176
rect 12433 4118 15903 4120
rect 12433 4115 12499 4118
rect 15837 4115 15903 4118
rect 2497 4042 2563 4045
rect 3509 4042 3575 4045
rect 2497 4040 3575 4042
rect 2497 3984 2502 4040
rect 2558 3984 3514 4040
rect 3570 3984 3575 4040
rect 2497 3982 3575 3984
rect 2497 3979 2563 3982
rect 3509 3979 3575 3982
rect 4061 4042 4127 4045
rect 16481 4042 16547 4045
rect 4061 4040 16547 4042
rect 4061 3984 4066 4040
rect 4122 3984 16486 4040
rect 16542 3984 16547 4040
rect 4061 3982 16547 3984
rect 4061 3979 4127 3982
rect 16481 3979 16547 3982
rect 2405 3906 2471 3909
rect 4981 3906 5047 3909
rect 2405 3904 5047 3906
rect 2405 3848 2410 3904
rect 2466 3848 4986 3904
rect 5042 3848 5047 3904
rect 2405 3846 5047 3848
rect 2405 3843 2471 3846
rect 4981 3843 5047 3846
rect 8201 3906 8267 3909
rect 12433 3906 12499 3909
rect 8201 3904 12499 3906
rect 8201 3848 8206 3904
rect 8262 3848 12438 3904
rect 12494 3848 12499 3904
rect 8201 3846 12499 3848
rect 8201 3843 8267 3846
rect 12433 3843 12499 3846
rect 12617 3906 12683 3909
rect 15285 3906 15351 3909
rect 12617 3904 15351 3906
rect 12617 3848 12622 3904
rect 12678 3848 15290 3904
rect 15346 3848 15351 3904
rect 12617 3846 15351 3848
rect 12617 3843 12683 3846
rect 15285 3843 15351 3846
rect 7562 3840 7878 3841
rect 7562 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7878 3840
rect 7562 3775 7878 3776
rect 2589 3770 2655 3773
rect 2454 3768 2655 3770
rect 2454 3712 2594 3768
rect 2650 3712 2655 3768
rect 2454 3710 2655 3712
rect 2454 3400 2514 3710
rect 2589 3707 2655 3710
rect 2773 3770 2839 3773
rect 4153 3770 4219 3773
rect 2773 3768 4219 3770
rect 2773 3712 2778 3768
rect 2834 3712 4158 3768
rect 4214 3712 4219 3768
rect 2773 3710 4219 3712
rect 2773 3707 2839 3710
rect 4153 3707 4219 3710
rect 9213 3770 9279 3773
rect 11789 3770 11855 3773
rect 9213 3768 11855 3770
rect 9213 3712 9218 3768
rect 9274 3712 11794 3768
rect 11850 3712 11855 3768
rect 9213 3710 11855 3712
rect 9213 3707 9279 3710
rect 11789 3707 11855 3710
rect 5533 3634 5599 3637
rect 15653 3634 15719 3637
rect 5533 3632 15719 3634
rect 5533 3576 5538 3632
rect 5594 3576 15658 3632
rect 15714 3576 15719 3632
rect 5533 3574 15719 3576
rect 5533 3571 5599 3574
rect 15653 3571 15719 3574
rect 2865 3498 2931 3501
rect 5533 3498 5599 3501
rect 2865 3496 5599 3498
rect 2865 3440 2870 3496
rect 2926 3440 5538 3496
rect 5594 3440 5599 3496
rect 2865 3438 5599 3440
rect 2865 3435 2931 3438
rect 5533 3435 5599 3438
rect 6913 3498 6979 3501
rect 15193 3498 15259 3501
rect 6913 3496 15259 3498
rect 6913 3440 6918 3496
rect 6974 3440 15198 3496
rect 15254 3440 15259 3496
rect 6913 3438 15259 3440
rect 6913 3435 6979 3438
rect 15193 3435 15259 3438
rect 9213 3362 9279 3365
rect 13353 3362 13419 3365
rect 9213 3360 13419 3362
rect 9213 3304 9218 3360
rect 9274 3304 13358 3360
rect 13414 3304 13419 3360
rect 9213 3302 13419 3304
rect 9213 3299 9279 3302
rect 13353 3299 13419 3302
rect 3562 3296 3878 3297
rect 3562 3232 3568 3296
rect 3632 3232 3648 3296
rect 3712 3232 3728 3296
rect 3792 3232 3808 3296
rect 3872 3232 3878 3296
rect 3562 3231 3878 3232
rect 8562 3296 8878 3297
rect 8562 3232 8568 3296
rect 8632 3232 8648 3296
rect 8712 3232 8728 3296
rect 8792 3232 8808 3296
rect 8872 3232 8878 3296
rect 8562 3231 8878 3232
rect 13537 3226 13603 3229
rect 9078 3224 13603 3226
rect 9078 3168 13542 3224
rect 13598 3168 13603 3224
rect 9078 3166 13603 3168
rect 2405 3090 2471 3093
rect 3509 3090 3575 3093
rect 2405 3088 3575 3090
rect 2405 3032 2410 3088
rect 2466 3032 3514 3088
rect 3570 3032 3575 3088
rect 2405 3030 3575 3032
rect 2405 3027 2471 3030
rect 3509 3027 3575 3030
rect 5901 3090 5967 3093
rect 9078 3090 9138 3166
rect 13537 3163 13603 3166
rect 5901 3088 9138 3090
rect 5901 3032 5906 3088
rect 5962 3032 9138 3088
rect 5901 3030 9138 3032
rect 9213 3090 9279 3093
rect 10133 3090 10199 3093
rect 9213 3088 10199 3090
rect 9213 3032 9218 3088
rect 9274 3032 10138 3088
rect 10194 3032 10199 3088
rect 9213 3030 10199 3032
rect 5901 3027 5967 3030
rect 9213 3027 9279 3030
rect 10133 3027 10199 3030
rect 3325 2954 3391 2957
rect 8109 2954 8175 2957
rect 3325 2952 8175 2954
rect 3325 2896 3330 2952
rect 3386 2896 8114 2952
rect 8170 2896 8175 2952
rect 3325 2894 8175 2896
rect 3325 2891 3391 2894
rect 8109 2891 8175 2894
rect 9622 2892 9628 2956
rect 9692 2954 9698 2956
rect 12341 2954 12407 2957
rect 9692 2952 12407 2954
rect 9692 2896 12346 2952
rect 12402 2896 12407 2952
rect 9692 2894 12407 2896
rect 9692 2892 9698 2894
rect 12341 2891 12407 2894
rect 12525 2954 12591 2957
rect 12893 2954 12959 2957
rect 12525 2952 12959 2954
rect 12525 2896 12530 2952
rect 12586 2896 12898 2952
rect 12954 2896 12959 2952
rect 12525 2894 12959 2896
rect 12525 2891 12591 2894
rect 12893 2891 12959 2894
rect 7281 2818 7347 2821
rect 12249 2818 12315 2821
rect 12801 2818 12867 2821
rect 6870 2816 7347 2818
rect 6870 2760 7286 2816
rect 7342 2760 7347 2816
rect 6870 2758 7347 2760
rect 4061 2682 4127 2685
rect 6870 2682 6930 2758
rect 7281 2755 7347 2758
rect 9262 2816 12315 2818
rect 9262 2760 12254 2816
rect 12310 2760 12315 2816
rect 9262 2758 12315 2760
rect 7562 2752 7878 2753
rect 7562 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7878 2752
rect 7562 2687 7878 2688
rect 4061 2680 6930 2682
rect 4061 2624 4066 2680
rect 4122 2624 6930 2680
rect 4061 2622 6930 2624
rect 8017 2682 8083 2685
rect 9262 2682 9322 2758
rect 12249 2755 12315 2758
rect 12390 2816 12867 2818
rect 12390 2760 12806 2816
rect 12862 2760 12867 2816
rect 12390 2758 12867 2760
rect 8017 2680 9322 2682
rect 8017 2624 8022 2680
rect 8078 2624 9322 2680
rect 8017 2622 9322 2624
rect 9397 2682 9463 2685
rect 12390 2682 12450 2758
rect 12801 2755 12867 2758
rect 9397 2680 12450 2682
rect 9397 2624 9402 2680
rect 9458 2624 12450 2680
rect 9397 2622 12450 2624
rect 14549 2682 14615 2685
rect 14549 2680 16866 2682
rect 14549 2624 14554 2680
rect 14610 2624 16866 2680
rect 14549 2622 16866 2624
rect 4061 2619 4127 2622
rect 8017 2619 8083 2622
rect 9397 2619 9463 2622
rect 14549 2619 14615 2622
rect 6913 2546 6979 2549
rect 14457 2546 14523 2549
rect 6913 2544 14523 2546
rect 6913 2488 6918 2544
rect 6974 2488 14462 2544
rect 14518 2488 14523 2544
rect 6913 2486 14523 2488
rect 6913 2483 6979 2486
rect 14457 2483 14523 2486
rect 6729 2410 6795 2413
rect 6729 2408 12450 2410
rect 6729 2352 6734 2408
rect 6790 2352 12450 2408
rect 6729 2350 12450 2352
rect 6729 2347 6795 2350
rect 12390 2274 12450 2350
rect 16021 2274 16087 2277
rect 12390 2272 16087 2274
rect 12390 2216 16026 2272
rect 16082 2216 16087 2272
rect 12390 2214 16087 2216
rect 16021 2211 16087 2214
rect 3562 2208 3878 2209
rect 3562 2144 3568 2208
rect 3632 2144 3648 2208
rect 3712 2144 3728 2208
rect 3792 2144 3808 2208
rect 3872 2144 3878 2208
rect 3562 2143 3878 2144
rect 8562 2208 8878 2209
rect 8562 2144 8568 2208
rect 8632 2144 8648 2208
rect 8712 2144 8728 2208
rect 8792 2144 8808 2208
rect 8872 2144 8878 2208
rect 8562 2143 8878 2144
rect 5625 2138 5691 2141
rect 8385 2138 8451 2141
rect 5625 2136 8451 2138
rect 5625 2080 5630 2136
rect 5686 2080 8390 2136
rect 8446 2080 8451 2136
rect 5625 2078 8451 2080
rect 5625 2075 5691 2078
rect 8385 2075 8451 2078
rect 9029 2138 9095 2141
rect 12157 2138 12223 2141
rect 9029 2136 12223 2138
rect 9029 2080 9034 2136
rect 9090 2080 12162 2136
rect 12218 2080 12223 2136
rect 9029 2078 12223 2080
rect 9029 2075 9095 2078
rect 12157 2075 12223 2078
rect 6085 2002 6151 2005
rect 9622 2002 9628 2004
rect 6085 2000 9628 2002
rect 6085 1944 6090 2000
rect 6146 1944 9628 2000
rect 6085 1942 9628 1944
rect 6085 1939 6151 1942
rect 9622 1940 9628 1942
rect 9692 1940 9698 2004
rect 4245 1866 4311 1869
rect 14549 1866 14615 1869
rect 4245 1864 14615 1866
rect 4245 1808 4250 1864
rect 4306 1808 14554 1864
rect 14610 1808 14615 1864
rect 4245 1806 14615 1808
rect 4245 1803 4311 1806
rect 14549 1803 14615 1806
rect 10593 1730 10659 1733
rect 8710 1728 10659 1730
rect 8710 1672 10598 1728
rect 10654 1672 10659 1728
rect 8710 1670 10659 1672
rect 7562 1664 7878 1665
rect 7562 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7878 1664
rect 7562 1599 7878 1600
rect 473 1594 539 1597
rect 1853 1594 1919 1597
rect 473 1592 1919 1594
rect 473 1536 478 1592
rect 534 1536 1858 1592
rect 1914 1536 1919 1592
rect 473 1534 1919 1536
rect 473 1531 539 1534
rect 1853 1531 1919 1534
rect 2313 1594 2379 1597
rect 4521 1594 4587 1597
rect 2313 1592 4587 1594
rect 2313 1536 2318 1592
rect 2374 1536 4526 1592
rect 4582 1536 4587 1592
rect 2313 1534 4587 1536
rect 2313 1531 2379 1534
rect 4521 1531 4587 1534
rect 1025 1458 1091 1461
rect 3141 1458 3207 1461
rect 1025 1456 3207 1458
rect 1025 1400 1030 1456
rect 1086 1400 3146 1456
rect 3202 1400 3207 1456
rect 1025 1398 3207 1400
rect 1025 1395 1091 1398
rect 3141 1395 3207 1398
rect 6269 1458 6335 1461
rect 8710 1458 8770 1670
rect 10593 1667 10659 1670
rect 14457 1730 14523 1733
rect 16665 1730 16731 1733
rect 14457 1728 16731 1730
rect 14457 1672 14462 1728
rect 14518 1672 16670 1728
rect 16726 1672 16731 1728
rect 14457 1670 16731 1672
rect 14457 1667 14523 1670
rect 16665 1667 16731 1670
rect 9213 1594 9279 1597
rect 16573 1594 16639 1597
rect 9213 1592 16639 1594
rect 9213 1536 9218 1592
rect 9274 1536 16578 1592
rect 16634 1536 16639 1592
rect 9213 1534 16639 1536
rect 9213 1531 9279 1534
rect 16573 1531 16639 1534
rect 6269 1456 8770 1458
rect 6269 1400 6274 1456
rect 6330 1400 8770 1456
rect 6269 1398 8770 1400
rect 8937 1458 9003 1461
rect 11881 1458 11947 1461
rect 8937 1456 11947 1458
rect 8937 1400 8942 1456
rect 8998 1400 11886 1456
rect 11942 1400 11947 1456
rect 8937 1398 11947 1400
rect 6269 1395 6335 1398
rect 8937 1395 9003 1398
rect 11881 1395 11947 1398
rect 16665 1458 16731 1461
rect 16806 1458 16866 2622
rect 16665 1456 16866 1458
rect 16665 1400 16670 1456
rect 16726 1400 16866 1456
rect 16665 1398 16866 1400
rect 16665 1395 16731 1398
rect 1117 1322 1183 1325
rect 4245 1322 4311 1325
rect 1117 1320 4311 1322
rect 1117 1264 1122 1320
rect 1178 1264 4250 1320
rect 4306 1264 4311 1320
rect 1117 1262 4311 1264
rect 1117 1259 1183 1262
rect 4245 1259 4311 1262
rect 7373 1322 7439 1325
rect 11329 1322 11395 1325
rect 7373 1320 11395 1322
rect 7373 1264 7378 1320
rect 7434 1264 11334 1320
rect 11390 1264 11395 1320
rect 7373 1262 11395 1264
rect 7373 1259 7439 1262
rect 11329 1259 11395 1262
rect 841 1186 907 1189
rect 2957 1186 3023 1189
rect 841 1184 3023 1186
rect 841 1128 846 1184
rect 902 1128 2962 1184
rect 3018 1128 3023 1184
rect 841 1126 3023 1128
rect 841 1123 907 1126
rect 2957 1123 3023 1126
rect 9121 1186 9187 1189
rect 12985 1186 13051 1189
rect 9121 1184 13051 1186
rect 9121 1128 9126 1184
rect 9182 1128 12990 1184
rect 13046 1128 13051 1184
rect 9121 1126 13051 1128
rect 9121 1123 9187 1126
rect 12985 1123 13051 1126
rect 3562 1120 3878 1121
rect 3562 1056 3568 1120
rect 3632 1056 3648 1120
rect 3712 1056 3728 1120
rect 3792 1056 3808 1120
rect 3872 1056 3878 1120
rect 3562 1055 3878 1056
rect 8562 1120 8878 1121
rect 8562 1056 8568 1120
rect 8632 1056 8648 1120
rect 8712 1056 8728 1120
rect 8792 1056 8808 1120
rect 8872 1056 8878 1120
rect 8562 1055 8878 1056
rect 4797 914 4863 917
rect 16113 914 16179 917
rect 4797 912 16179 914
rect 4797 856 4802 912
rect 4858 856 16118 912
rect 16174 856 16179 912
rect 4797 854 16179 856
rect 4797 851 4863 854
rect 16113 851 16179 854
rect 289 778 355 781
rect 6729 778 6795 781
rect 289 776 6795 778
rect 289 720 294 776
rect 350 720 6734 776
rect 6790 720 6795 776
rect 289 718 6795 720
rect 289 715 355 718
rect 6729 715 6795 718
rect 8385 778 8451 781
rect 10317 778 10383 781
rect 8385 776 10383 778
rect 8385 720 8390 776
rect 8446 720 10322 776
rect 10378 720 10383 776
rect 8385 718 10383 720
rect 8385 715 8451 718
rect 10317 715 10383 718
rect 4981 642 5047 645
rect 16389 642 16455 645
rect 4981 640 16455 642
rect 4981 584 4986 640
rect 5042 584 16394 640
rect 16450 584 16455 640
rect 4981 582 16455 584
rect 4981 579 5047 582
rect 16389 579 16455 582
rect 6545 506 6611 509
rect 12617 506 12683 509
rect 6545 504 12683 506
rect 6545 448 6550 504
rect 6606 448 12622 504
rect 12678 448 12683 504
rect 6545 446 12683 448
rect 6545 443 6611 446
rect 12617 443 12683 446
rect 4061 370 4127 373
rect 14273 370 14339 373
rect 4061 368 14339 370
rect 4061 312 4066 368
rect 4122 312 14278 368
rect 14334 312 14339 368
rect 4061 310 14339 312
rect 4061 307 4127 310
rect 14273 307 14339 310
rect 6085 98 6151 101
rect 16297 98 16363 101
rect 6085 96 16363 98
rect 6085 40 6090 96
rect 6146 40 16302 96
rect 16358 40 16363 96
rect 6085 38 16363 40
rect 6085 35 6151 38
rect 16297 35 16363 38
<< via3 >>
rect 2568 15804 2632 15808
rect 2568 15748 2572 15804
rect 2572 15748 2628 15804
rect 2628 15748 2632 15804
rect 2568 15744 2632 15748
rect 2648 15804 2712 15808
rect 2648 15748 2652 15804
rect 2652 15748 2708 15804
rect 2708 15748 2712 15804
rect 2648 15744 2712 15748
rect 2728 15804 2792 15808
rect 2728 15748 2732 15804
rect 2732 15748 2788 15804
rect 2788 15748 2792 15804
rect 2728 15744 2792 15748
rect 2808 15804 2872 15808
rect 2808 15748 2812 15804
rect 2812 15748 2868 15804
rect 2868 15748 2872 15804
rect 2808 15744 2872 15748
rect 7568 15804 7632 15808
rect 7568 15748 7572 15804
rect 7572 15748 7628 15804
rect 7628 15748 7632 15804
rect 7568 15744 7632 15748
rect 7648 15804 7712 15808
rect 7648 15748 7652 15804
rect 7652 15748 7708 15804
rect 7708 15748 7712 15804
rect 7648 15744 7712 15748
rect 7728 15804 7792 15808
rect 7728 15748 7732 15804
rect 7732 15748 7788 15804
rect 7788 15748 7792 15804
rect 7728 15744 7792 15748
rect 7808 15804 7872 15808
rect 7808 15748 7812 15804
rect 7812 15748 7868 15804
rect 7868 15748 7872 15804
rect 7808 15744 7872 15748
rect 3568 15260 3632 15264
rect 3568 15204 3572 15260
rect 3572 15204 3628 15260
rect 3628 15204 3632 15260
rect 3568 15200 3632 15204
rect 3648 15260 3712 15264
rect 3648 15204 3652 15260
rect 3652 15204 3708 15260
rect 3708 15204 3712 15260
rect 3648 15200 3712 15204
rect 3728 15260 3792 15264
rect 3728 15204 3732 15260
rect 3732 15204 3788 15260
rect 3788 15204 3792 15260
rect 3728 15200 3792 15204
rect 3808 15260 3872 15264
rect 3808 15204 3812 15260
rect 3812 15204 3868 15260
rect 3868 15204 3872 15260
rect 3808 15200 3872 15204
rect 8568 15260 8632 15264
rect 8568 15204 8572 15260
rect 8572 15204 8628 15260
rect 8628 15204 8632 15260
rect 8568 15200 8632 15204
rect 8648 15260 8712 15264
rect 8648 15204 8652 15260
rect 8652 15204 8708 15260
rect 8708 15204 8712 15260
rect 8648 15200 8712 15204
rect 8728 15260 8792 15264
rect 8728 15204 8732 15260
rect 8732 15204 8788 15260
rect 8788 15204 8792 15260
rect 8728 15200 8792 15204
rect 8808 15260 8872 15264
rect 8808 15204 8812 15260
rect 8812 15204 8868 15260
rect 8868 15204 8872 15260
rect 8808 15200 8872 15204
rect 2568 14716 2632 14720
rect 2568 14660 2572 14716
rect 2572 14660 2628 14716
rect 2628 14660 2632 14716
rect 2568 14656 2632 14660
rect 2648 14716 2712 14720
rect 2648 14660 2652 14716
rect 2652 14660 2708 14716
rect 2708 14660 2712 14716
rect 2648 14656 2712 14660
rect 2728 14716 2792 14720
rect 2728 14660 2732 14716
rect 2732 14660 2788 14716
rect 2788 14660 2792 14716
rect 2728 14656 2792 14660
rect 2808 14716 2872 14720
rect 2808 14660 2812 14716
rect 2812 14660 2868 14716
rect 2868 14660 2872 14716
rect 2808 14656 2872 14660
rect 7568 14716 7632 14720
rect 7568 14660 7572 14716
rect 7572 14660 7628 14716
rect 7628 14660 7632 14716
rect 7568 14656 7632 14660
rect 7648 14716 7712 14720
rect 7648 14660 7652 14716
rect 7652 14660 7708 14716
rect 7708 14660 7712 14716
rect 7648 14656 7712 14660
rect 7728 14716 7792 14720
rect 7728 14660 7732 14716
rect 7732 14660 7788 14716
rect 7788 14660 7792 14716
rect 7728 14656 7792 14660
rect 7808 14716 7872 14720
rect 7808 14660 7812 14716
rect 7812 14660 7868 14716
rect 7868 14660 7872 14716
rect 7808 14656 7872 14660
rect 3568 14172 3632 14176
rect 3568 14116 3572 14172
rect 3572 14116 3628 14172
rect 3628 14116 3632 14172
rect 3568 14112 3632 14116
rect 3648 14172 3712 14176
rect 3648 14116 3652 14172
rect 3652 14116 3708 14172
rect 3708 14116 3712 14172
rect 3648 14112 3712 14116
rect 3728 14172 3792 14176
rect 3728 14116 3732 14172
rect 3732 14116 3788 14172
rect 3788 14116 3792 14172
rect 3728 14112 3792 14116
rect 3808 14172 3872 14176
rect 3808 14116 3812 14172
rect 3812 14116 3868 14172
rect 3868 14116 3872 14172
rect 3808 14112 3872 14116
rect 8568 14172 8632 14176
rect 8568 14116 8572 14172
rect 8572 14116 8628 14172
rect 8628 14116 8632 14172
rect 8568 14112 8632 14116
rect 8648 14172 8712 14176
rect 8648 14116 8652 14172
rect 8652 14116 8708 14172
rect 8708 14116 8712 14172
rect 8648 14112 8712 14116
rect 8728 14172 8792 14176
rect 8728 14116 8732 14172
rect 8732 14116 8788 14172
rect 8788 14116 8792 14172
rect 8728 14112 8792 14116
rect 8808 14172 8872 14176
rect 8808 14116 8812 14172
rect 8812 14116 8868 14172
rect 8868 14116 8872 14172
rect 8808 14112 8872 14116
rect 2568 13628 2632 13632
rect 2568 13572 2572 13628
rect 2572 13572 2628 13628
rect 2628 13572 2632 13628
rect 2568 13568 2632 13572
rect 2648 13628 2712 13632
rect 2648 13572 2652 13628
rect 2652 13572 2708 13628
rect 2708 13572 2712 13628
rect 2648 13568 2712 13572
rect 2728 13628 2792 13632
rect 2728 13572 2732 13628
rect 2732 13572 2788 13628
rect 2788 13572 2792 13628
rect 2728 13568 2792 13572
rect 2808 13628 2872 13632
rect 2808 13572 2812 13628
rect 2812 13572 2868 13628
rect 2868 13572 2872 13628
rect 2808 13568 2872 13572
rect 7568 13628 7632 13632
rect 7568 13572 7572 13628
rect 7572 13572 7628 13628
rect 7628 13572 7632 13628
rect 7568 13568 7632 13572
rect 7648 13628 7712 13632
rect 7648 13572 7652 13628
rect 7652 13572 7708 13628
rect 7708 13572 7712 13628
rect 7648 13568 7712 13572
rect 7728 13628 7792 13632
rect 7728 13572 7732 13628
rect 7732 13572 7788 13628
rect 7788 13572 7792 13628
rect 7728 13568 7792 13572
rect 7808 13628 7872 13632
rect 7808 13572 7812 13628
rect 7812 13572 7868 13628
rect 7868 13572 7872 13628
rect 7808 13568 7872 13572
rect 3568 13084 3632 13088
rect 3568 13028 3572 13084
rect 3572 13028 3628 13084
rect 3628 13028 3632 13084
rect 3568 13024 3632 13028
rect 3648 13084 3712 13088
rect 3648 13028 3652 13084
rect 3652 13028 3708 13084
rect 3708 13028 3712 13084
rect 3648 13024 3712 13028
rect 3728 13084 3792 13088
rect 3728 13028 3732 13084
rect 3732 13028 3788 13084
rect 3788 13028 3792 13084
rect 3728 13024 3792 13028
rect 3808 13084 3872 13088
rect 3808 13028 3812 13084
rect 3812 13028 3868 13084
rect 3868 13028 3872 13084
rect 3808 13024 3872 13028
rect 8568 13084 8632 13088
rect 8568 13028 8572 13084
rect 8572 13028 8628 13084
rect 8628 13028 8632 13084
rect 8568 13024 8632 13028
rect 8648 13084 8712 13088
rect 8648 13028 8652 13084
rect 8652 13028 8708 13084
rect 8708 13028 8712 13084
rect 8648 13024 8712 13028
rect 8728 13084 8792 13088
rect 8728 13028 8732 13084
rect 8732 13028 8788 13084
rect 8788 13028 8792 13084
rect 8728 13024 8792 13028
rect 8808 13084 8872 13088
rect 8808 13028 8812 13084
rect 8812 13028 8868 13084
rect 8868 13028 8872 13084
rect 8808 13024 8872 13028
rect 2268 12684 2332 12748
rect 2568 12540 2632 12544
rect 2568 12484 2572 12540
rect 2572 12484 2628 12540
rect 2628 12484 2632 12540
rect 2568 12480 2632 12484
rect 2648 12540 2712 12544
rect 2648 12484 2652 12540
rect 2652 12484 2708 12540
rect 2708 12484 2712 12540
rect 2648 12480 2712 12484
rect 2728 12540 2792 12544
rect 2728 12484 2732 12540
rect 2732 12484 2788 12540
rect 2788 12484 2792 12540
rect 2728 12480 2792 12484
rect 2808 12540 2872 12544
rect 2808 12484 2812 12540
rect 2812 12484 2868 12540
rect 2868 12484 2872 12540
rect 2808 12480 2872 12484
rect 7568 12540 7632 12544
rect 7568 12484 7572 12540
rect 7572 12484 7628 12540
rect 7628 12484 7632 12540
rect 7568 12480 7632 12484
rect 7648 12540 7712 12544
rect 7648 12484 7652 12540
rect 7652 12484 7708 12540
rect 7708 12484 7712 12540
rect 7648 12480 7712 12484
rect 7728 12540 7792 12544
rect 7728 12484 7732 12540
rect 7732 12484 7788 12540
rect 7788 12484 7792 12540
rect 7728 12480 7792 12484
rect 7808 12540 7872 12544
rect 7808 12484 7812 12540
rect 7812 12484 7868 12540
rect 7868 12484 7872 12540
rect 7808 12480 7872 12484
rect 9260 12004 9324 12068
rect 3568 11996 3632 12000
rect 3568 11940 3572 11996
rect 3572 11940 3628 11996
rect 3628 11940 3632 11996
rect 3568 11936 3632 11940
rect 3648 11996 3712 12000
rect 3648 11940 3652 11996
rect 3652 11940 3708 11996
rect 3708 11940 3712 11996
rect 3648 11936 3712 11940
rect 3728 11996 3792 12000
rect 3728 11940 3732 11996
rect 3732 11940 3788 11996
rect 3788 11940 3792 11996
rect 3728 11936 3792 11940
rect 3808 11996 3872 12000
rect 3808 11940 3812 11996
rect 3812 11940 3868 11996
rect 3868 11940 3872 11996
rect 3808 11936 3872 11940
rect 8568 11996 8632 12000
rect 8568 11940 8572 11996
rect 8572 11940 8628 11996
rect 8628 11940 8632 11996
rect 8568 11936 8632 11940
rect 8648 11996 8712 12000
rect 8648 11940 8652 11996
rect 8652 11940 8708 11996
rect 8708 11940 8712 11996
rect 8648 11936 8712 11940
rect 8728 11996 8792 12000
rect 8728 11940 8732 11996
rect 8732 11940 8788 11996
rect 8788 11940 8792 11996
rect 8728 11936 8792 11940
rect 8808 11996 8872 12000
rect 8808 11940 8812 11996
rect 8812 11940 8868 11996
rect 8868 11940 8872 11996
rect 8808 11936 8872 11940
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 7568 11452 7632 11456
rect 7568 11396 7572 11452
rect 7572 11396 7628 11452
rect 7628 11396 7632 11452
rect 7568 11392 7632 11396
rect 7648 11452 7712 11456
rect 7648 11396 7652 11452
rect 7652 11396 7708 11452
rect 7708 11396 7712 11452
rect 7648 11392 7712 11396
rect 7728 11452 7792 11456
rect 7728 11396 7732 11452
rect 7732 11396 7788 11452
rect 7788 11396 7792 11452
rect 7728 11392 7792 11396
rect 7808 11452 7872 11456
rect 7808 11396 7812 11452
rect 7812 11396 7868 11452
rect 7868 11396 7872 11452
rect 7808 11392 7872 11396
rect 3568 10908 3632 10912
rect 3568 10852 3572 10908
rect 3572 10852 3628 10908
rect 3628 10852 3632 10908
rect 3568 10848 3632 10852
rect 3648 10908 3712 10912
rect 3648 10852 3652 10908
rect 3652 10852 3708 10908
rect 3708 10852 3712 10908
rect 3648 10848 3712 10852
rect 3728 10908 3792 10912
rect 3728 10852 3732 10908
rect 3732 10852 3788 10908
rect 3788 10852 3792 10908
rect 3728 10848 3792 10852
rect 3808 10908 3872 10912
rect 3808 10852 3812 10908
rect 3812 10852 3868 10908
rect 3868 10852 3872 10908
rect 3808 10848 3872 10852
rect 8568 10908 8632 10912
rect 8568 10852 8572 10908
rect 8572 10852 8628 10908
rect 8628 10852 8632 10908
rect 8568 10848 8632 10852
rect 8648 10908 8712 10912
rect 8648 10852 8652 10908
rect 8652 10852 8708 10908
rect 8708 10852 8712 10908
rect 8648 10848 8712 10852
rect 8728 10908 8792 10912
rect 8728 10852 8732 10908
rect 8732 10852 8788 10908
rect 8788 10852 8792 10908
rect 8728 10848 8792 10852
rect 8808 10908 8872 10912
rect 8808 10852 8812 10908
rect 8812 10852 8868 10908
rect 8868 10852 8872 10908
rect 8808 10848 8872 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 7568 10364 7632 10368
rect 7568 10308 7572 10364
rect 7572 10308 7628 10364
rect 7628 10308 7632 10364
rect 7568 10304 7632 10308
rect 7648 10364 7712 10368
rect 7648 10308 7652 10364
rect 7652 10308 7708 10364
rect 7708 10308 7712 10364
rect 7648 10304 7712 10308
rect 7728 10364 7792 10368
rect 7728 10308 7732 10364
rect 7732 10308 7788 10364
rect 7788 10308 7792 10364
rect 7728 10304 7792 10308
rect 7808 10364 7872 10368
rect 7808 10308 7812 10364
rect 7812 10308 7868 10364
rect 7868 10308 7872 10364
rect 7808 10304 7872 10308
rect 3568 9820 3632 9824
rect 3568 9764 3572 9820
rect 3572 9764 3628 9820
rect 3628 9764 3632 9820
rect 3568 9760 3632 9764
rect 3648 9820 3712 9824
rect 3648 9764 3652 9820
rect 3652 9764 3708 9820
rect 3708 9764 3712 9820
rect 3648 9760 3712 9764
rect 3728 9820 3792 9824
rect 3728 9764 3732 9820
rect 3732 9764 3788 9820
rect 3788 9764 3792 9820
rect 3728 9760 3792 9764
rect 3808 9820 3872 9824
rect 3808 9764 3812 9820
rect 3812 9764 3868 9820
rect 3868 9764 3872 9820
rect 3808 9760 3872 9764
rect 8568 9820 8632 9824
rect 8568 9764 8572 9820
rect 8572 9764 8628 9820
rect 8628 9764 8632 9820
rect 8568 9760 8632 9764
rect 8648 9820 8712 9824
rect 8648 9764 8652 9820
rect 8652 9764 8708 9820
rect 8708 9764 8712 9820
rect 8648 9760 8712 9764
rect 8728 9820 8792 9824
rect 8728 9764 8732 9820
rect 8732 9764 8788 9820
rect 8788 9764 8792 9820
rect 8728 9760 8792 9764
rect 8808 9820 8872 9824
rect 8808 9764 8812 9820
rect 8812 9764 8868 9820
rect 8868 9764 8872 9820
rect 8808 9760 8872 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 7568 9276 7632 9280
rect 7568 9220 7572 9276
rect 7572 9220 7628 9276
rect 7628 9220 7632 9276
rect 7568 9216 7632 9220
rect 7648 9276 7712 9280
rect 7648 9220 7652 9276
rect 7652 9220 7708 9276
rect 7708 9220 7712 9276
rect 7648 9216 7712 9220
rect 7728 9276 7792 9280
rect 7728 9220 7732 9276
rect 7732 9220 7788 9276
rect 7788 9220 7792 9276
rect 7728 9216 7792 9220
rect 7808 9276 7872 9280
rect 7808 9220 7812 9276
rect 7812 9220 7868 9276
rect 7868 9220 7872 9276
rect 7808 9216 7872 9220
rect 3568 8732 3632 8736
rect 3568 8676 3572 8732
rect 3572 8676 3628 8732
rect 3628 8676 3632 8732
rect 3568 8672 3632 8676
rect 3648 8732 3712 8736
rect 3648 8676 3652 8732
rect 3652 8676 3708 8732
rect 3708 8676 3712 8732
rect 3648 8672 3712 8676
rect 3728 8732 3792 8736
rect 3728 8676 3732 8732
rect 3732 8676 3788 8732
rect 3788 8676 3792 8732
rect 3728 8672 3792 8676
rect 3808 8732 3872 8736
rect 3808 8676 3812 8732
rect 3812 8676 3868 8732
rect 3868 8676 3872 8732
rect 3808 8672 3872 8676
rect 8568 8732 8632 8736
rect 8568 8676 8572 8732
rect 8572 8676 8628 8732
rect 8628 8676 8632 8732
rect 8568 8672 8632 8676
rect 8648 8732 8712 8736
rect 8648 8676 8652 8732
rect 8652 8676 8708 8732
rect 8708 8676 8712 8732
rect 8648 8672 8712 8676
rect 8728 8732 8792 8736
rect 8728 8676 8732 8732
rect 8732 8676 8788 8732
rect 8788 8676 8792 8732
rect 8728 8672 8792 8676
rect 8808 8732 8872 8736
rect 8808 8676 8812 8732
rect 8812 8676 8868 8732
rect 8868 8676 8872 8732
rect 8808 8672 8872 8676
rect 6868 8196 6932 8260
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 7568 8188 7632 8192
rect 7568 8132 7572 8188
rect 7572 8132 7628 8188
rect 7628 8132 7632 8188
rect 7568 8128 7632 8132
rect 7648 8188 7712 8192
rect 7648 8132 7652 8188
rect 7652 8132 7708 8188
rect 7708 8132 7712 8188
rect 7648 8128 7712 8132
rect 7728 8188 7792 8192
rect 7728 8132 7732 8188
rect 7732 8132 7788 8188
rect 7788 8132 7792 8188
rect 7728 8128 7792 8132
rect 7808 8188 7872 8192
rect 7808 8132 7812 8188
rect 7812 8132 7868 8188
rect 7868 8132 7872 8188
rect 7808 8128 7872 8132
rect 2268 7924 2332 7988
rect 3568 7644 3632 7648
rect 3568 7588 3572 7644
rect 3572 7588 3628 7644
rect 3628 7588 3632 7644
rect 3568 7584 3632 7588
rect 3648 7644 3712 7648
rect 3648 7588 3652 7644
rect 3652 7588 3708 7644
rect 3708 7588 3712 7644
rect 3648 7584 3712 7588
rect 3728 7644 3792 7648
rect 3728 7588 3732 7644
rect 3732 7588 3788 7644
rect 3788 7588 3792 7644
rect 3728 7584 3792 7588
rect 3808 7644 3872 7648
rect 3808 7588 3812 7644
rect 3812 7588 3868 7644
rect 3868 7588 3872 7644
rect 3808 7584 3872 7588
rect 8568 7644 8632 7648
rect 8568 7588 8572 7644
rect 8572 7588 8628 7644
rect 8628 7588 8632 7644
rect 8568 7584 8632 7588
rect 8648 7644 8712 7648
rect 8648 7588 8652 7644
rect 8652 7588 8708 7644
rect 8708 7588 8712 7644
rect 8648 7584 8712 7588
rect 8728 7644 8792 7648
rect 8728 7588 8732 7644
rect 8732 7588 8788 7644
rect 8788 7588 8792 7644
rect 8728 7584 8792 7588
rect 8808 7644 8872 7648
rect 8808 7588 8812 7644
rect 8812 7588 8868 7644
rect 8868 7588 8872 7644
rect 8808 7584 8872 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 7568 7100 7632 7104
rect 7568 7044 7572 7100
rect 7572 7044 7628 7100
rect 7628 7044 7632 7100
rect 7568 7040 7632 7044
rect 7648 7100 7712 7104
rect 7648 7044 7652 7100
rect 7652 7044 7708 7100
rect 7708 7044 7712 7100
rect 7648 7040 7712 7044
rect 7728 7100 7792 7104
rect 7728 7044 7732 7100
rect 7732 7044 7788 7100
rect 7788 7044 7792 7100
rect 7728 7040 7792 7044
rect 7808 7100 7872 7104
rect 7808 7044 7812 7100
rect 7812 7044 7868 7100
rect 7868 7044 7872 7100
rect 7808 7040 7872 7044
rect 3568 6556 3632 6560
rect 3568 6500 3572 6556
rect 3572 6500 3628 6556
rect 3628 6500 3632 6556
rect 3568 6496 3632 6500
rect 3648 6556 3712 6560
rect 3648 6500 3652 6556
rect 3652 6500 3708 6556
rect 3708 6500 3712 6556
rect 3648 6496 3712 6500
rect 3728 6556 3792 6560
rect 3728 6500 3732 6556
rect 3732 6500 3788 6556
rect 3788 6500 3792 6556
rect 3728 6496 3792 6500
rect 3808 6556 3872 6560
rect 3808 6500 3812 6556
rect 3812 6500 3868 6556
rect 3868 6500 3872 6556
rect 3808 6496 3872 6500
rect 8568 6556 8632 6560
rect 8568 6500 8572 6556
rect 8572 6500 8628 6556
rect 8628 6500 8632 6556
rect 8568 6496 8632 6500
rect 8648 6556 8712 6560
rect 8648 6500 8652 6556
rect 8652 6500 8708 6556
rect 8708 6500 8712 6556
rect 8648 6496 8712 6500
rect 8728 6556 8792 6560
rect 8728 6500 8732 6556
rect 8732 6500 8788 6556
rect 8788 6500 8792 6556
rect 8728 6496 8792 6500
rect 8808 6556 8872 6560
rect 8808 6500 8812 6556
rect 8812 6500 8868 6556
rect 8868 6500 8872 6556
rect 8808 6496 8872 6500
rect 2268 6488 2332 6492
rect 2268 6432 2282 6488
rect 2282 6432 2332 6488
rect 2268 6428 2332 6432
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 7568 6012 7632 6016
rect 7568 5956 7572 6012
rect 7572 5956 7628 6012
rect 7628 5956 7632 6012
rect 7568 5952 7632 5956
rect 7648 6012 7712 6016
rect 7648 5956 7652 6012
rect 7652 5956 7708 6012
rect 7708 5956 7712 6012
rect 7648 5952 7712 5956
rect 7728 6012 7792 6016
rect 7728 5956 7732 6012
rect 7732 5956 7788 6012
rect 7788 5956 7792 6012
rect 7728 5952 7792 5956
rect 7808 6012 7872 6016
rect 7808 5956 7812 6012
rect 7812 5956 7868 6012
rect 7868 5956 7872 6012
rect 7808 5952 7872 5956
rect 6868 5476 6932 5540
rect 3568 5468 3632 5472
rect 3568 5412 3572 5468
rect 3572 5412 3628 5468
rect 3628 5412 3632 5468
rect 3568 5408 3632 5412
rect 3648 5468 3712 5472
rect 3648 5412 3652 5468
rect 3652 5412 3708 5468
rect 3708 5412 3712 5468
rect 3648 5408 3712 5412
rect 3728 5468 3792 5472
rect 3728 5412 3732 5468
rect 3732 5412 3788 5468
rect 3788 5412 3792 5468
rect 3728 5408 3792 5412
rect 3808 5468 3872 5472
rect 3808 5412 3812 5468
rect 3812 5412 3868 5468
rect 3868 5412 3872 5468
rect 3808 5408 3872 5412
rect 8568 5468 8632 5472
rect 8568 5412 8572 5468
rect 8572 5412 8628 5468
rect 8628 5412 8632 5468
rect 8568 5408 8632 5412
rect 8648 5468 8712 5472
rect 8648 5412 8652 5468
rect 8652 5412 8708 5468
rect 8708 5412 8712 5468
rect 8648 5408 8712 5412
rect 8728 5468 8792 5472
rect 8728 5412 8732 5468
rect 8732 5412 8788 5468
rect 8788 5412 8792 5468
rect 8728 5408 8792 5412
rect 8808 5468 8872 5472
rect 8808 5412 8812 5468
rect 8812 5412 8868 5468
rect 8868 5412 8872 5468
rect 8808 5408 8872 5412
rect 7568 4924 7632 4928
rect 7568 4868 7572 4924
rect 7572 4868 7628 4924
rect 7628 4868 7632 4924
rect 7568 4864 7632 4868
rect 7648 4924 7712 4928
rect 7648 4868 7652 4924
rect 7652 4868 7708 4924
rect 7708 4868 7712 4924
rect 7648 4864 7712 4868
rect 7728 4924 7792 4928
rect 7728 4868 7732 4924
rect 7732 4868 7788 4924
rect 7788 4868 7792 4924
rect 7728 4864 7792 4868
rect 7808 4924 7872 4928
rect 7808 4868 7812 4924
rect 7812 4868 7868 4924
rect 7868 4868 7872 4924
rect 7808 4864 7872 4868
rect 3568 4380 3632 4384
rect 3568 4324 3572 4380
rect 3572 4324 3628 4380
rect 3628 4324 3632 4380
rect 3568 4320 3632 4324
rect 3648 4380 3712 4384
rect 3648 4324 3652 4380
rect 3652 4324 3708 4380
rect 3708 4324 3712 4380
rect 3648 4320 3712 4324
rect 3728 4380 3792 4384
rect 3728 4324 3732 4380
rect 3732 4324 3788 4380
rect 3788 4324 3792 4380
rect 3728 4320 3792 4324
rect 3808 4380 3872 4384
rect 3808 4324 3812 4380
rect 3812 4324 3868 4380
rect 3868 4324 3872 4380
rect 3808 4320 3872 4324
rect 8568 4380 8632 4384
rect 8568 4324 8572 4380
rect 8572 4324 8628 4380
rect 8628 4324 8632 4380
rect 8568 4320 8632 4324
rect 8648 4380 8712 4384
rect 8648 4324 8652 4380
rect 8652 4324 8708 4380
rect 8708 4324 8712 4380
rect 8648 4320 8712 4324
rect 8728 4380 8792 4384
rect 8728 4324 8732 4380
rect 8732 4324 8788 4380
rect 8788 4324 8792 4380
rect 8728 4320 8792 4324
rect 8808 4380 8872 4384
rect 8808 4324 8812 4380
rect 8812 4324 8868 4380
rect 8868 4324 8872 4380
rect 8808 4320 8872 4324
rect 7568 3836 7632 3840
rect 7568 3780 7572 3836
rect 7572 3780 7628 3836
rect 7628 3780 7632 3836
rect 7568 3776 7632 3780
rect 7648 3836 7712 3840
rect 7648 3780 7652 3836
rect 7652 3780 7708 3836
rect 7708 3780 7712 3836
rect 7648 3776 7712 3780
rect 7728 3836 7792 3840
rect 7728 3780 7732 3836
rect 7732 3780 7788 3836
rect 7788 3780 7792 3836
rect 7728 3776 7792 3780
rect 7808 3836 7872 3840
rect 7808 3780 7812 3836
rect 7812 3780 7868 3836
rect 7868 3780 7872 3836
rect 7808 3776 7872 3780
rect 3568 3292 3632 3296
rect 3568 3236 3572 3292
rect 3572 3236 3628 3292
rect 3628 3236 3632 3292
rect 3568 3232 3632 3236
rect 3648 3292 3712 3296
rect 3648 3236 3652 3292
rect 3652 3236 3708 3292
rect 3708 3236 3712 3292
rect 3648 3232 3712 3236
rect 3728 3292 3792 3296
rect 3728 3236 3732 3292
rect 3732 3236 3788 3292
rect 3788 3236 3792 3292
rect 3728 3232 3792 3236
rect 3808 3292 3872 3296
rect 3808 3236 3812 3292
rect 3812 3236 3868 3292
rect 3868 3236 3872 3292
rect 3808 3232 3872 3236
rect 8568 3292 8632 3296
rect 8568 3236 8572 3292
rect 8572 3236 8628 3292
rect 8628 3236 8632 3292
rect 8568 3232 8632 3236
rect 8648 3292 8712 3296
rect 8648 3236 8652 3292
rect 8652 3236 8708 3292
rect 8708 3236 8712 3292
rect 8648 3232 8712 3236
rect 8728 3292 8792 3296
rect 8728 3236 8732 3292
rect 8732 3236 8788 3292
rect 8788 3236 8792 3292
rect 8728 3232 8792 3236
rect 8808 3292 8872 3296
rect 8808 3236 8812 3292
rect 8812 3236 8868 3292
rect 8868 3236 8872 3292
rect 8808 3232 8872 3236
rect 9628 2892 9692 2956
rect 7568 2748 7632 2752
rect 7568 2692 7572 2748
rect 7572 2692 7628 2748
rect 7628 2692 7632 2748
rect 7568 2688 7632 2692
rect 7648 2748 7712 2752
rect 7648 2692 7652 2748
rect 7652 2692 7708 2748
rect 7708 2692 7712 2748
rect 7648 2688 7712 2692
rect 7728 2748 7792 2752
rect 7728 2692 7732 2748
rect 7732 2692 7788 2748
rect 7788 2692 7792 2748
rect 7728 2688 7792 2692
rect 7808 2748 7872 2752
rect 7808 2692 7812 2748
rect 7812 2692 7868 2748
rect 7868 2692 7872 2748
rect 7808 2688 7872 2692
rect 3568 2204 3632 2208
rect 3568 2148 3572 2204
rect 3572 2148 3628 2204
rect 3628 2148 3632 2204
rect 3568 2144 3632 2148
rect 3648 2204 3712 2208
rect 3648 2148 3652 2204
rect 3652 2148 3708 2204
rect 3708 2148 3712 2204
rect 3648 2144 3712 2148
rect 3728 2204 3792 2208
rect 3728 2148 3732 2204
rect 3732 2148 3788 2204
rect 3788 2148 3792 2204
rect 3728 2144 3792 2148
rect 3808 2204 3872 2208
rect 3808 2148 3812 2204
rect 3812 2148 3868 2204
rect 3868 2148 3872 2204
rect 3808 2144 3872 2148
rect 8568 2204 8632 2208
rect 8568 2148 8572 2204
rect 8572 2148 8628 2204
rect 8628 2148 8632 2204
rect 8568 2144 8632 2148
rect 8648 2204 8712 2208
rect 8648 2148 8652 2204
rect 8652 2148 8708 2204
rect 8708 2148 8712 2204
rect 8648 2144 8712 2148
rect 8728 2204 8792 2208
rect 8728 2148 8732 2204
rect 8732 2148 8788 2204
rect 8788 2148 8792 2204
rect 8728 2144 8792 2148
rect 8808 2204 8872 2208
rect 8808 2148 8812 2204
rect 8812 2148 8868 2204
rect 8868 2148 8872 2204
rect 8808 2144 8872 2148
rect 9628 1940 9692 2004
rect 7568 1660 7632 1664
rect 7568 1604 7572 1660
rect 7572 1604 7628 1660
rect 7628 1604 7632 1660
rect 7568 1600 7632 1604
rect 7648 1660 7712 1664
rect 7648 1604 7652 1660
rect 7652 1604 7708 1660
rect 7708 1604 7712 1660
rect 7648 1600 7712 1604
rect 7728 1660 7792 1664
rect 7728 1604 7732 1660
rect 7732 1604 7788 1660
rect 7788 1604 7792 1660
rect 7728 1600 7792 1604
rect 7808 1660 7872 1664
rect 7808 1604 7812 1660
rect 7812 1604 7868 1660
rect 7868 1604 7872 1660
rect 7808 1600 7872 1604
rect 3568 1116 3632 1120
rect 3568 1060 3572 1116
rect 3572 1060 3628 1116
rect 3628 1060 3632 1116
rect 3568 1056 3632 1060
rect 3648 1116 3712 1120
rect 3648 1060 3652 1116
rect 3652 1060 3708 1116
rect 3708 1060 3712 1116
rect 3648 1056 3712 1060
rect 3728 1116 3792 1120
rect 3728 1060 3732 1116
rect 3732 1060 3788 1116
rect 3788 1060 3792 1116
rect 3728 1056 3792 1060
rect 3808 1116 3872 1120
rect 3808 1060 3812 1116
rect 3812 1060 3868 1116
rect 3868 1060 3872 1116
rect 3808 1056 3872 1060
rect 8568 1116 8632 1120
rect 8568 1060 8572 1116
rect 8572 1060 8628 1116
rect 8628 1060 8632 1116
rect 8568 1056 8632 1060
rect 8648 1116 8712 1120
rect 8648 1060 8652 1116
rect 8652 1060 8708 1116
rect 8708 1060 8712 1116
rect 8648 1056 8712 1060
rect 8728 1116 8792 1120
rect 8728 1060 8732 1116
rect 8732 1060 8788 1116
rect 8788 1060 8792 1116
rect 8728 1056 8792 1060
rect 8808 1116 8872 1120
rect 8808 1060 8812 1116
rect 8812 1060 8868 1116
rect 8868 1060 8872 1116
rect 8808 1056 8872 1060
<< metal4 >>
rect 2560 15808 2880 15824
rect 2560 15744 2568 15808
rect 2632 15744 2648 15808
rect 2712 15744 2728 15808
rect 2792 15744 2808 15808
rect 2872 15744 2880 15808
rect 2560 14720 2880 15744
rect 2560 14656 2568 14720
rect 2632 14656 2648 14720
rect 2712 14656 2728 14720
rect 2792 14656 2808 14720
rect 2872 14656 2880 14720
rect 2560 13632 2880 14656
rect 2560 13568 2568 13632
rect 2632 13568 2648 13632
rect 2712 13568 2728 13632
rect 2792 13568 2808 13632
rect 2872 13568 2880 13632
rect 2560 13206 2880 13568
rect 2560 12970 2602 13206
rect 2838 12970 2880 13206
rect 2267 12748 2333 12749
rect 2267 12684 2268 12748
rect 2332 12684 2333 12748
rect 2267 12683 2333 12684
rect 2270 12018 2330 12683
rect 2560 12544 2880 12970
rect 2560 12480 2568 12544
rect 2632 12480 2648 12544
rect 2712 12480 2728 12544
rect 2792 12480 2808 12544
rect 2872 12480 2880 12544
rect 2560 11456 2880 12480
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9206 2880 9216
rect 2560 8970 2602 9206
rect 2838 8970 2880 9206
rect 2560 8192 2880 8970
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2267 7988 2333 7989
rect 2267 7924 2268 7988
rect 2332 7924 2333 7988
rect 2267 7923 2333 7924
rect 2270 6493 2330 7923
rect 2560 7104 2880 8128
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2267 6492 2333 6493
rect 2267 6428 2268 6492
rect 2332 6428 2333 6492
rect 2267 6427 2333 6428
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5206 2880 5952
rect 2560 4970 2602 5206
rect 2838 4970 2880 5206
rect 2560 4893 2880 4970
rect 3560 15264 3880 15824
rect 3560 15200 3568 15264
rect 3632 15200 3648 15264
rect 3712 15200 3728 15264
rect 3792 15200 3808 15264
rect 3872 15200 3880 15264
rect 3560 14206 3880 15200
rect 3560 14176 3602 14206
rect 3838 14176 3880 14206
rect 3560 14112 3568 14176
rect 3872 14112 3880 14176
rect 3560 13970 3602 14112
rect 3838 13970 3880 14112
rect 3560 13088 3880 13970
rect 3560 13024 3568 13088
rect 3632 13024 3648 13088
rect 3712 13024 3728 13088
rect 3792 13024 3808 13088
rect 3872 13024 3880 13088
rect 3560 12000 3880 13024
rect 3560 11936 3568 12000
rect 3632 11936 3648 12000
rect 3712 11936 3728 12000
rect 3792 11936 3808 12000
rect 3872 11936 3880 12000
rect 3560 10912 3880 11936
rect 3560 10848 3568 10912
rect 3632 10848 3648 10912
rect 3712 10848 3728 10912
rect 3792 10848 3808 10912
rect 3872 10848 3880 10912
rect 3560 10206 3880 10848
rect 3560 9970 3602 10206
rect 3838 9970 3880 10206
rect 3560 9824 3880 9970
rect 3560 9760 3568 9824
rect 3632 9760 3648 9824
rect 3712 9760 3728 9824
rect 3792 9760 3808 9824
rect 3872 9760 3880 9824
rect 3560 8736 3880 9760
rect 3560 8672 3568 8736
rect 3632 8672 3648 8736
rect 3712 8672 3728 8736
rect 3792 8672 3808 8736
rect 3872 8672 3880 8736
rect 3560 7648 3880 8672
rect 3560 7584 3568 7648
rect 3632 7584 3648 7648
rect 3712 7584 3728 7648
rect 3792 7584 3808 7648
rect 3872 7584 3880 7648
rect 3560 6560 3880 7584
rect 3560 6496 3568 6560
rect 3632 6496 3648 6560
rect 3712 6496 3728 6560
rect 3792 6496 3808 6560
rect 3872 6496 3880 6560
rect 3560 6206 3880 6496
rect 3560 5970 3602 6206
rect 3838 5970 3880 6206
rect 3560 5472 3880 5970
rect 3560 5408 3568 5472
rect 3632 5408 3648 5472
rect 3712 5408 3728 5472
rect 3792 5408 3808 5472
rect 3872 5408 3880 5472
rect 3560 4384 3880 5408
rect 3560 4320 3568 4384
rect 3632 4320 3648 4384
rect 3712 4320 3728 4384
rect 3792 4320 3808 4384
rect 3872 4320 3880 4384
rect 1996 4206 2276 4248
rect 1996 3970 2018 4206
rect 2254 3970 2276 4206
rect 1996 3928 2276 3970
rect 3560 3296 3880 4320
rect 1256 3206 1536 3248
rect 1256 2970 1278 3206
rect 1514 2970 1536 3206
rect 1256 2928 1536 2970
rect 3560 3232 3568 3296
rect 3632 3232 3648 3296
rect 3712 3232 3728 3296
rect 3792 3232 3808 3296
rect 3872 3232 3880 3296
rect 3560 2208 3880 3232
rect 3560 2144 3568 2208
rect 3632 2206 3648 2208
rect 3712 2206 3728 2208
rect 3792 2206 3808 2208
rect 3872 2144 3880 2208
rect 3560 1970 3602 2144
rect 3838 1970 3880 2144
rect 3560 1120 3880 1970
rect 3560 1056 3568 1120
rect 3632 1056 3648 1120
rect 3712 1056 3728 1120
rect 3792 1056 3808 1120
rect 3872 1056 3880 1120
rect 3560 1040 3880 1056
rect 4560 3206 4880 15824
rect 4560 2970 4602 3206
rect 4838 2970 4880 3206
rect 4560 1040 4880 2970
rect 5560 4206 5880 15824
rect 7560 15808 7880 15824
rect 7560 15744 7568 15808
rect 7632 15744 7648 15808
rect 7712 15744 7728 15808
rect 7792 15744 7808 15808
rect 7872 15744 7880 15808
rect 7560 14720 7880 15744
rect 7560 14656 7568 14720
rect 7632 14656 7648 14720
rect 7712 14656 7728 14720
rect 7792 14656 7808 14720
rect 7872 14656 7880 14720
rect 7560 13632 7880 14656
rect 7560 13568 7568 13632
rect 7632 13568 7648 13632
rect 7712 13568 7728 13632
rect 7792 13568 7808 13632
rect 7872 13568 7880 13632
rect 7560 13206 7880 13568
rect 7560 12970 7602 13206
rect 7838 12970 7880 13206
rect 7560 12544 7880 12970
rect 7560 12480 7568 12544
rect 7632 12480 7648 12544
rect 7712 12480 7728 12544
rect 7792 12480 7808 12544
rect 7872 12480 7880 12544
rect 7560 11456 7880 12480
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 7560 10368 7880 11392
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 9280 7880 10304
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 9206 7880 9216
rect 7560 8970 7602 9206
rect 7838 8970 7880 9206
rect 6867 8260 6933 8261
rect 6867 8196 6868 8260
rect 6932 8196 6933 8260
rect 6867 8195 6933 8196
rect 6870 5541 6930 8195
rect 7560 8192 7880 8970
rect 7560 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7880 8192
rect 7560 7104 7880 8128
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 6016 7880 7040
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 6867 5540 6933 5541
rect 6867 5476 6868 5540
rect 6932 5476 6933 5540
rect 6867 5475 6933 5476
rect 5560 3970 5602 4206
rect 5838 3970 5880 4206
rect 5560 1040 5880 3970
rect 7560 5206 7880 5952
rect 7560 4970 7602 5206
rect 7838 4970 7880 5206
rect 7560 4928 7880 4970
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 7560 3840 7880 4864
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 2752 7880 3776
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 1664 7880 2688
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 7560 1206 7880 1600
rect 7560 970 7602 1206
rect 7838 970 7880 1206
rect 8560 15264 8880 15824
rect 8560 15200 8568 15264
rect 8632 15200 8648 15264
rect 8712 15200 8728 15264
rect 8792 15200 8808 15264
rect 8872 15200 8880 15264
rect 8560 14206 8880 15200
rect 8560 14176 8602 14206
rect 8838 14176 8880 14206
rect 8560 14112 8568 14176
rect 8872 14112 8880 14176
rect 8560 13970 8602 14112
rect 8838 13970 8880 14112
rect 8560 13088 8880 13970
rect 8560 13024 8568 13088
rect 8632 13024 8648 13088
rect 8712 13024 8728 13088
rect 8792 13024 8808 13088
rect 8872 13024 8880 13088
rect 8560 12000 8880 13024
rect 9259 12068 9325 12069
rect 9259 12018 9260 12068
rect 9324 12018 9325 12068
rect 8560 11936 8568 12000
rect 8632 11936 8648 12000
rect 8712 11936 8728 12000
rect 8792 11936 8808 12000
rect 8872 11936 8880 12000
rect 8560 10912 8880 11936
rect 8560 10848 8568 10912
rect 8632 10848 8648 10912
rect 8712 10848 8728 10912
rect 8792 10848 8808 10912
rect 8872 10848 8880 10912
rect 8560 10206 8880 10848
rect 8560 9970 8602 10206
rect 8838 9970 8880 10206
rect 8560 9824 8880 9970
rect 8560 9760 8568 9824
rect 8632 9760 8648 9824
rect 8712 9760 8728 9824
rect 8792 9760 8808 9824
rect 8872 9760 8880 9824
rect 8560 8736 8880 9760
rect 8560 8672 8568 8736
rect 8632 8672 8648 8736
rect 8712 8672 8728 8736
rect 8792 8672 8808 8736
rect 8872 8672 8880 8736
rect 8560 7648 8880 8672
rect 8560 7584 8568 7648
rect 8632 7584 8648 7648
rect 8712 7584 8728 7648
rect 8792 7584 8808 7648
rect 8872 7584 8880 7648
rect 8560 6560 8880 7584
rect 8560 6496 8568 6560
rect 8632 6496 8648 6560
rect 8712 6496 8728 6560
rect 8792 6496 8808 6560
rect 8872 6496 8880 6560
rect 8560 6206 8880 6496
rect 8560 5970 8602 6206
rect 8838 5970 8880 6206
rect 8560 5472 8880 5970
rect 8560 5408 8568 5472
rect 8632 5408 8648 5472
rect 8712 5408 8728 5472
rect 8792 5408 8808 5472
rect 8872 5408 8880 5472
rect 8560 4384 8880 5408
rect 8560 4320 8568 4384
rect 8632 4320 8648 4384
rect 8712 4320 8728 4384
rect 8792 4320 8808 4384
rect 8872 4320 8880 4384
rect 8560 3296 8880 4320
rect 8560 3232 8568 3296
rect 8632 3232 8648 3296
rect 8712 3232 8728 3296
rect 8792 3232 8808 3296
rect 8872 3232 8880 3296
rect 8560 2208 8880 3232
rect 9627 2956 9693 2957
rect 9627 2892 9628 2956
rect 9692 2892 9693 2956
rect 9627 2891 9693 2892
rect 8560 2144 8568 2208
rect 8632 2206 8648 2208
rect 8712 2206 8728 2208
rect 8792 2206 8808 2208
rect 8872 2144 8880 2208
rect 8560 1970 8602 2144
rect 8838 1970 8880 2144
rect 9630 2005 9690 2891
rect 8560 1120 8880 1970
rect 9627 2004 9693 2005
rect 9627 1940 9628 2004
rect 9692 1940 9693 2004
rect 9627 1939 9693 1940
rect 8560 1056 8568 1120
rect 8632 1056 8648 1120
rect 8712 1056 8728 1120
rect 8792 1056 8808 1120
rect 8872 1056 8880 1120
rect 8560 1040 8880 1056
rect 7560 928 7880 970
<< via4 >>
rect 2602 12970 2838 13206
rect 2182 11782 2418 12018
rect 2602 8970 2838 9206
rect 2602 4970 2838 5206
rect 3602 14176 3838 14206
rect 3602 14112 3632 14176
rect 3632 14112 3648 14176
rect 3648 14112 3712 14176
rect 3712 14112 3728 14176
rect 3728 14112 3792 14176
rect 3792 14112 3808 14176
rect 3808 14112 3838 14176
rect 3602 13970 3838 14112
rect 3602 9970 3838 10206
rect 3602 5970 3838 6206
rect 2018 3970 2254 4206
rect 1278 2970 1514 3206
rect 3602 2144 3632 2206
rect 3632 2144 3648 2206
rect 3648 2144 3712 2206
rect 3712 2144 3728 2206
rect 3728 2144 3792 2206
rect 3792 2144 3808 2206
rect 3808 2144 3838 2206
rect 3602 1970 3838 2144
rect 4602 2970 4838 3206
rect 7602 12970 7838 13206
rect 7602 8970 7838 9206
rect 5602 3970 5838 4206
rect 7602 4970 7838 5206
rect 7602 970 7838 1206
rect 8602 14176 8838 14206
rect 8602 14112 8632 14176
rect 8632 14112 8648 14176
rect 8648 14112 8712 14176
rect 8712 14112 8728 14176
rect 8728 14112 8792 14176
rect 8792 14112 8808 14176
rect 8808 14112 8838 14176
rect 8602 13970 8838 14112
rect 9174 12004 9260 12018
rect 9260 12004 9324 12018
rect 9324 12004 9410 12018
rect 9174 11782 9410 12004
rect 8602 9970 8838 10206
rect 8602 5970 8838 6206
rect 8602 2144 8632 2206
rect 8632 2144 8648 2206
rect 8648 2144 8712 2206
rect 8712 2144 8728 2206
rect 8728 2144 8792 2206
rect 8792 2144 8808 2206
rect 8808 2144 8838 2206
rect 8602 1970 8838 2144
<< metal5 >>
rect 872 14206 9892 14248
rect 872 13970 3602 14206
rect 3838 13970 8602 14206
rect 8838 13970 9892 14206
rect 872 13928 9892 13970
rect 872 13206 9892 13248
rect 872 12970 2602 13206
rect 2838 12970 7602 13206
rect 7838 12970 9892 13206
rect 872 12928 9892 12970
rect 2140 12018 9452 12060
rect 2140 11782 2182 12018
rect 2418 11782 9174 12018
rect 9410 11782 9452 12018
rect 2140 11740 9452 11782
rect 872 10206 9892 10248
rect 872 9970 3602 10206
rect 3838 9970 8602 10206
rect 8838 9970 9892 10206
rect 872 9928 9892 9970
rect 872 9206 9892 9248
rect 872 8970 2602 9206
rect 2838 8970 7602 9206
rect 7838 8970 9892 9206
rect 872 8928 9892 8970
rect 872 6206 9892 6248
rect 872 5970 3602 6206
rect 3838 5970 8602 6206
rect 8838 5970 9892 6206
rect 872 5928 9892 5970
rect 872 5206 9892 5248
rect 872 4970 2602 5206
rect 2838 4970 7602 5206
rect 7838 4970 9892 5206
rect 872 4928 9892 4970
rect 872 4206 9892 4248
rect 872 3970 2018 4206
rect 2254 3970 5602 4206
rect 5838 3970 9892 4206
rect 872 3928 9892 3970
rect 872 3206 9892 3248
rect 872 2970 1278 3206
rect 1514 2970 4602 3206
rect 4838 2970 9892 3206
rect 872 2928 9892 2970
rect 872 2206 9892 2248
rect 872 1970 3602 2206
rect 3838 1970 8602 2206
rect 8838 1970 9892 2206
rect 872 1928 9892 1970
rect 872 1206 9892 1248
rect 872 970 7602 1206
rect 7838 970 9892 1206
rect 872 928 9892 970
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 3312 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 3772 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1663720911
transform 1 0 4416 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 5060 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52
timestamp 1663720911
transform 1 0 5704 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1663720911
transform 1 0 6164 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64
timestamp 1663720911
transform 1 0 6808 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 7452 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80
timestamp 1663720911
transform 1 0 8280 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1663720911
transform 1 0 9200 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1663720911
transform 1 0 3312 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_31
timestamp 1663720911
transform 1 0 3772 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1663720911
transform 1 0 4416 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1663720911
transform 1 0 5060 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1663720911
transform 1 0 5704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_59
timestamp 1663720911
transform 1 0 6348 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_66 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 6992 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1663720911
transform 1 0 8096 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_80
timestamp 1663720911
transform 1 0 8280 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 1663720911
transform 1 0 8740 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1663720911
transform 1 0 9384 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1663720911
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_31
timestamp 1663720911
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_38
timestamp 1663720911
transform 1 0 4416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_45
timestamp 1663720911
transform 1 0 5060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_52
timestamp 1663720911
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1663720911
transform 1 0 6164 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_64
timestamp 1663720911
transform 1 0 6808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_76
timestamp 1663720911
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_80
timestamp 1663720911
transform 1 0 8280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_84
timestamp 1663720911
transform 1 0 8648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_91 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1663720911
transform 1 0 3312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_31
timestamp 1663720911
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_38
timestamp 1663720911
transform 1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_42
timestamp 1663720911
transform 1 0 4784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_46
timestamp 1663720911
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_53
timestamp 1663720911
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_60
timestamp 1663720911
transform 1 0 6440 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_67
timestamp 1663720911
transform 1 0 7084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_73
timestamp 1663720911
transform 1 0 7636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1663720911
transform 1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_80
timestamp 1663720911
transform 1 0 8280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1663720911
transform 1 0 9384 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1663720911
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_31
timestamp 1663720911
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_38
timestamp 1663720911
transform 1 0 4416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_45
timestamp 1663720911
transform 1 0 5060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_52
timestamp 1663720911
transform 1 0 5704 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_57
timestamp 1663720911
transform 1 0 6164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_66
timestamp 1663720911
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_73
timestamp 1663720911
transform 1 0 7636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_80
timestamp 1663720911
transform 1 0 8280 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_92
timestamp 1663720911
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_26
timestamp 1663720911
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1663720911
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1663720911
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1663720911
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_59
timestamp 1663720911
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_66
timestamp 1663720911
transform 1 0 6992 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_72
timestamp 1663720911
transform 1 0 7544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_76
timestamp 1663720911
transform 1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_80
timestamp 1663720911
transform 1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1663720911
transform 1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1663720911
transform 1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_31
timestamp 1663720911
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_35
timestamp 1663720911
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_45
timestamp 1663720911
transform 1 0 5060 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_52
timestamp 1663720911
transform 1 0 5704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1663720911
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_65
timestamp 1663720911
transform 1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_72
timestamp 1663720911
transform 1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_84
timestamp 1663720911
transform 1 0 8648 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_92
timestamp 1663720911
transform 1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_26
timestamp 1663720911
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_30
timestamp 1663720911
transform 1 0 3680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1663720911
transform 1 0 4048 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1663720911
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_53
timestamp 1663720911
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_65
timestamp 1663720911
transform 1 0 6900 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1663720911
transform 1 0 7728 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_78
timestamp 1663720911
transform 1 0 8096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_80
timestamp 1663720911
transform 1 0 8280 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_86
timestamp 1663720911
transform 1 0 8832 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_91
timestamp 1663720911
transform 1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1663720911
transform 1 0 1196 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1663720911
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_12
timestamp 1663720911
transform 1 0 2024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_16
timestamp 1663720911
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1663720911
transform 1 0 3036 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1663720911
transform 1 0 3404 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1663720911
transform 1 0 3588 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1663720911
transform 1 0 5612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_55
timestamp 1663720911
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_57
timestamp 1663720911
transform 1 0 6164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_63
timestamp 1663720911
transform 1 0 6716 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1663720911
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1663720911
transform 1 0 8740 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_91
timestamp 1663720911
transform 1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1663720911
transform 1 0 1196 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_9
timestamp 1663720911
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_17
timestamp 1663720911
transform 1 0 2484 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_25
timestamp 1663720911
transform 1 0 3220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_46
timestamp 1663720911
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1663720911
transform 1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1663720911
transform 1 0 6164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_61
timestamp 1663720911
transform 1 0 6532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_88
timestamp 1663720911
transform 1 0 9016 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1663720911
transform 1 0 1196 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1663720911
transform 1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1663720911
transform 1 0 3588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_52
timestamp 1663720911
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1663720911
transform 1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1663720911
transform 1 0 8740 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_92
timestamp 1663720911
transform 1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1663720911
transform 1 0 1196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1663720911
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1663720911
transform 1 0 3680 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1663720911
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1663720911
transform 1 0 6164 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1663720911
transform 1 0 8740 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1663720911
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1663720911
transform 1 0 1196 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1663720911
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1663720911
transform 1 0 3588 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_39
timestamp 1663720911
transform 1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_67
timestamp 1663720911
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1663720911
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1663720911
transform 1 0 8556 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1663720911
transform 1 0 8740 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_92
timestamp 1663720911
transform 1 0 9384 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1663720911
transform 1 0 1196 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1663720911
transform 1 0 1564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_12
timestamp 1663720911
transform 1 0 2024 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_46
timestamp 1663720911
transform 1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1663720911
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1663720911
transform 1 0 6164 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_67
timestamp 1663720911
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp 1663720911
transform 1 0 9384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1663720911
transform 1 0 1196 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1663720911
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1663720911
transform 1 0 3588 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp 1663720911
transform 1 0 3956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_42
timestamp 1663720911
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1663720911
transform 1 0 5152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_67
timestamp 1663720911
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1663720911
transform 1 0 8004 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1663720911
transform 1 0 8556 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1663720911
transform 1 0 8740 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_91
timestamp 1663720911
transform 1 0 9292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1663720911
transform 1 0 1196 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_12
timestamp 1663720911
transform 1 0 2024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1663720911
transform 1 0 3128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1663720911
transform 1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1663720911
transform 1 0 6164 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 1663720911
transform 1 0 6992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_90
timestamp 1663720911
transform 1 0 9200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1663720911
transform 1 0 1196 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_12
timestamp 1663720911
transform 1 0 2024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1663720911
transform 1 0 3128 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1663720911
transform 1 0 3588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_51
timestamp 1663720911
transform 1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1663720911
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1663720911
transform 1 0 8740 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_92
timestamp 1663720911
transform 1 0 9384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1663720911
transform 1 0 1196 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1663720911
transform 1 0 1564 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1663720911
transform 1 0 2116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_43
timestamp 1663720911
transform 1 0 4876 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1663720911
transform 1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1663720911
transform 1 0 6164 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1663720911
transform 1 0 8740 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_92
timestamp 1663720911
transform 1 0 9384 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1663720911
transform 1 0 1196 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1663720911
transform 1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1663720911
transform 1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1663720911
transform 1 0 3588 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_45
timestamp 1663720911
transform 1 0 5060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_69
timestamp 1663720911
transform 1 0 7268 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_77
timestamp 1663720911
transform 1 0 8004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1663720911
transform 1 0 8464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1663720911
transform 1 0 8740 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_91
timestamp 1663720911
transform 1 0 9292 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1663720911
transform 1 0 1196 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 1663720911
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_30
timestamp 1663720911
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1663720911
transform 1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1663720911
transform 1 0 6164 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_79
timestamp 1663720911
transform 1 0 8188 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_91
timestamp 1663720911
transform 1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1663720911
transform 1 0 1196 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1663720911
transform 1 0 3312 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1663720911
transform 1 0 3588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 1663720911
transform 1 0 4048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_64
timestamp 1663720911
transform 1 0 6808 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_70
timestamp 1663720911
transform 1 0 7360 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1663720911
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1663720911
transform 1 0 8556 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1663720911
transform 1 0 8740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_92
timestamp 1663720911
transform 1 0 9384 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1663720911
transform 1 0 1196 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_13
timestamp 1663720911
transform 1 0 2116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_43
timestamp 1663720911
transform 1 0 4876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_47
timestamp 1663720911
transform 1 0 5244 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1663720911
transform 1 0 5888 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1663720911
transform 1 0 6164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_81
timestamp 1663720911
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_85
timestamp 1663720911
transform 1 0 8740 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp 1663720911
transform 1 0 9384 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1663720911
transform 1 0 1196 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1663720911
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1663720911
transform 1 0 3588 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_40
timestamp 1663720911
transform 1 0 4600 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_72
timestamp 1663720911
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_76
timestamp 1663720911
transform 1 0 7912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1663720911
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1663720911
transform 1 0 8740 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_91
timestamp 1663720911
transform 1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1663720911
transform 1 0 1196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_14
timestamp 1663720911
transform 1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_44
timestamp 1663720911
transform 1 0 4968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1663720911
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1663720911
transform 1 0 6164 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1663720911
transform 1 0 6532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_88
timestamp 1663720911
transform 1 0 9016 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1663720911
transform 1 0 1196 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1663720911
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_29
timestamp 1663720911
transform 1 0 3588 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_43
timestamp 1663720911
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_67
timestamp 1663720911
transform 1 0 7084 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1663720911
transform 1 0 8188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1663720911
transform 1 0 8556 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1663720911
transform 1 0 8740 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_92
timestamp 1663720911
transform 1 0 9384 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1663720911
transform 1 0 1196 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_8
timestamp 1663720911
transform 1 0 1656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_17
timestamp 1663720911
transform 1 0 2484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_26
timestamp 1663720911
transform 1 0 3312 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_38
timestamp 1663720911
transform 1 0 4416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1663720911
transform 1 0 5520 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1663720911
transform 1 0 6164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_61
timestamp 1663720911
transform 1 0 6532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_82
timestamp 1663720911
transform 1 0 8464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_92
timestamp 1663720911
transform 1 0 9384 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1663720911
transform 1 0 1196 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_10
timestamp 1663720911
transform 1 0 1840 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_18
timestamp 1663720911
transform 1 0 2576 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1663720911
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1663720911
transform 1 0 3588 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1663720911
transform 1 0 4692 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_54
timestamp 1663720911
transform 1 0 5888 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_57
timestamp 1663720911
transform 1 0 6164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 1663720911
transform 1 0 6532 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1663720911
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1663720911
transform 1 0 8740 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_91
timestamp 1663720911
transform 1 0 9292 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1663720911
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1663720911
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1663720911
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1663720911
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1663720911
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1663720911
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1663720911
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1663720911
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1663720911
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1663720911
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1663720911
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1663720911
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1663720911
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1663720911
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1663720911
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1663720911
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1663720911
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1663720911
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1663720911
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1663720911
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1663720911
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1663720911
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1663720911
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1663720911
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1663720911
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1663720911
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1663720911
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1663720911
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1663720911
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1663720911
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1663720911
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1663720911
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1663720911
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1663720911
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1663720911
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1663720911
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1663720911
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1663720911
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1663720911
transform 1 0 920 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1663720911
transform -1 0 9844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1663720911
transform 1 0 920 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1663720911
transform -1 0 9844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1663720911
transform 1 0 920 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1663720911
transform -1 0 9844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1663720911
transform 1 0 920 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1663720911
transform -1 0 9844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1663720911
transform 1 0 920 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1663720911
transform -1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1663720911
transform 1 0 920 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1663720911
transform -1 0 9844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1663720911
transform 1 0 920 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1663720911
transform -1 0 9844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1663720911
transform 1 0 920 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1663720911
transform -1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1663720911
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1663720911
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1663720911
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1663720911
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1663720911
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1663720911
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1663720911
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1663720911
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1663720911
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1663720911
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1663720911
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1663720911
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1663720911
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1663720911
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1663720911
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1663720911
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1663720911
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1663720911
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1663720911
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1663720911
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1663720911
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1663720911
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1663720911
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1663720911
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1663720911
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1663720911
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1663720911
transform 1 0 6072 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1663720911
transform 1 0 3496 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1663720911
transform 1 0 8648 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1663720911
transform 1 0 6072 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1663720911
transform 1 0 3496 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1663720911
transform 1 0 8648 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1663720911
transform 1 0 6072 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1663720911
transform 1 0 3496 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1663720911
transform 1 0 8648 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1663720911
transform 1 0 6072 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1663720911
transform 1 0 3496 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1663720911
transform 1 0 6072 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1663720911
transform 1 0 8648 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 6440 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 9384 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 8740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _090_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 3496 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1663720911
transform -1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _093_
timestamp 1663720911
transform 1 0 3496 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 9016 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 8096 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1663720911
transform -1 0 8740 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _097_
timestamp 1663720911
transform -1 0 8648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _098_
timestamp 1663720911
transform -1 0 9292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _099_
timestamp 1663720911
transform -1 0 6992 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _100_
timestamp 1663720911
transform 1 0 7176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1663720911
transform -1 0 9384 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 2024 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 6532 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 5336 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _106__5
timestamp 1663720911
transform -1 0 4416 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp 1663720911
transform -1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _108_
timestamp 1663720911
transform 1 0 7452 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _109_
timestamp 1663720911
transform 1 0 4784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _110_
timestamp 1663720911
transform 1 0 1564 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1663720911
transform -1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112__6
timestamp 1663720911
transform -1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _113_
timestamp 1663720911
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _114_
timestamp 1663720911
transform 1 0 5336 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1663720911
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116__7
timestamp 1663720911
transform -1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _117_
timestamp 1663720911
transform 1 0 4784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _118_
timestamp 1663720911
transform 1 0 8924 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1663720911
transform -1 0 6164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120__8
timestamp 1663720911
transform 1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _121_
timestamp 1663720911
transform 1 0 4784 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 1663720911
transform -1 0 2116 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1663720911
transform -1 0 3772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124__9
timestamp 1663720911
transform 1 0 4140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _125_
timestamp 1663720911
transform 1 0 4784 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _126_
timestamp 1663720911
transform 1 0 1564 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1663720911
transform -1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _128__10
timestamp 1663720911
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _129_
timestamp 1663720911
transform 1 0 4140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _130_
timestamp 1663720911
transform 1 0 2852 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1663720911
transform 1 0 6164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _132__11
timestamp 1663720911
transform 1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _133_
timestamp 1663720911
transform 1 0 5888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _134_
timestamp 1663720911
transform 1 0 5428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1663720911
transform 1 0 9108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136__12
timestamp 1663720911
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _137_
timestamp 1663720911
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _138_
timestamp 1663720911
transform 1 0 8924 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1663720911
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _140__13
timestamp 1663720911
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _141_
timestamp 1663720911
transform -1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _142_
timestamp 1663720911
transform -1 0 3312 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1663720911
transform -1 0 6348 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144__14
timestamp 1663720911
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _145_
timestamp 1663720911
transform 1 0 5428 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _146_
timestamp 1663720911
transform 1 0 8924 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1663720911
transform -1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148__1
timestamp 1663720911
transform -1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _149_
timestamp 1663720911
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _150_
timestamp 1663720911
transform 1 0 8924 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1663720911
transform 1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _152__2
timestamp 1663720911
transform -1 0 6900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _153_
timestamp 1663720911
transform -1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _154_
timestamp 1663720911
transform 1 0 7268 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1663720911
transform -1 0 8004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156__3
timestamp 1663720911
transform 1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _157_
timestamp 1663720911
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _158__4
timestamp 1663720911
transform 1 0 4140 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 2576 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _160_
timestamp 1663720911
transform 1 0 2484 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _161_
timestamp 1663720911
transform 1 0 4416 0 1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _162_
timestamp 1663720911
transform 1 0 5152 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _163_
timestamp 1663720911
transform 1 0 2760 0 -1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _164_
timestamp 1663720911
transform 1 0 3496 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _165_
timestamp 1663720911
transform 1 0 2484 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _166_
timestamp 1663720911
transform 1 0 5980 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _167_
timestamp 1663720911
transform 1 0 6348 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _168_
timestamp 1663720911
transform 1 0 6624 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _169_
timestamp 1663720911
transform 1 0 6348 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _170_
timestamp 1663720911
transform 1 0 6072 0 1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _171_
timestamp 1663720911
transform 1 0 6624 0 -1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__dfrtp_1  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 8464 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _173_
timestamp 1663720911
transform -1 0 3312 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _174_
timestamp 1663720911
transform -1 0 3312 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _175_
timestamp 1663720911
transform 1 0 1472 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _176_
timestamp 1663720911
transform 1 0 1472 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _177_
timestamp 1663720911
transform 1 0 3772 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _178_
timestamp 1663720911
transform -1 0 5704 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _179_
timestamp 1663720911
transform 1 0 4048 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _180_
timestamp 1663720911
transform -1 0 5152 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _181_
timestamp 1663720911
transform -1 0 3680 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _182_
timestamp 1663720911
transform 1 0 3772 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _183_
timestamp 1663720911
transform 1 0 6348 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _184_
timestamp 1663720911
transform 1 0 6532 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _185_
timestamp 1663720911
transform -1 0 8464 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 1663720911
transform 1 0 9016 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 1840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _188_
timestamp 1663720911
transform -1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_8  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 9384 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 5888 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock
timestamp 1663720911
transform -1 0 7268 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 1663720911
transform -1 0 9200 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__068_
timestamp 1663720911
transform -1 0 3312 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_clock
timestamp 1663720911
transform -1 0 3680 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_load
timestamp 1663720911
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__068_
timestamp 1663720911
transform 1 0 1472 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_clock
timestamp 1663720911
transform 1 0 5244 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_load
timestamp 1663720911
transform -1 0 7084 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 9200 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1663720911
transform -1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 9384 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 6808 0 1 5440
box -38 -48 1694 592
use gpio_logic_high  gpio_logic_high
timestamp 0
transform 1 0 1196 0 1 1680
box -1196 -1680 32804 15320
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1663720911
transform -1 0 8188 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1663720911
transform -1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1663720911
transform 1 0 2392 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1663720911
transform 1 0 1472 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1663720911
transform -1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1663720911
transform -1 0 8188 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1663720911
transform 1 0 4048 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1663720911
transform 1 0 1472 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1663720911
transform 1 0 2576 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1663720911
transform 1 0 6164 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1663720911
transform 1 0 5060 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1663720911
transform -1 0 8188 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1663720911
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1663720911
transform 1 0 3680 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1663720911
transform 1 0 3956 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1663720911
transform -1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1663720911
transform -1 0 5060 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1663720911
transform 1 0 2392 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output1
timestamp 1663720911
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 1663720911
transform -1 0 8648 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1663720911
transform 1 0 9016 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1663720911
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1663720911
transform 1 0 5520 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1663720911
transform 1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1663720911
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1663720911
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1663720911
transform 1 0 9016 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1663720911
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1663720911
transform -1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1663720911
transform 1 0 8004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1663720911
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1663720911
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  output15
timestamp 1663720911
transform 1 0 3588 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output16
timestamp 1663720911
transform -1 0 5888 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output17
timestamp 1663720911
transform 1 0 4232 0 1 4352
box -38 -48 866 592
<< labels >>
flabel metal2 s 938 16200 994 17000 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 0 nsew signal input
flabel metal2 s 5538 16200 5594 17000 0 FreeSans 224 90 0 0 gpio_defaults[10]
port 1 nsew signal input
flabel metal2 s 5998 16200 6054 17000 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 2 nsew signal input
flabel metal2 s 6458 16200 6514 17000 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 3 nsew signal input
flabel metal2 s 1398 16200 1454 17000 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 4 nsew signal input
flabel metal2 s 1858 16200 1914 17000 0 FreeSans 224 90 0 0 gpio_defaults[2]
port 5 nsew signal input
flabel metal2 s 2318 16200 2374 17000 0 FreeSans 224 90 0 0 gpio_defaults[3]
port 6 nsew signal input
flabel metal2 s 2778 16200 2834 17000 0 FreeSans 224 90 0 0 gpio_defaults[4]
port 7 nsew signal input
flabel metal2 s 3238 16200 3294 17000 0 FreeSans 224 90 0 0 gpio_defaults[5]
port 8 nsew signal input
flabel metal2 s 3698 16200 3754 17000 0 FreeSans 224 90 0 0 gpio_defaults[6]
port 9 nsew signal input
flabel metal2 s 4158 16200 4214 17000 0 FreeSans 224 90 0 0 gpio_defaults[7]
port 10 nsew signal input
flabel metal2 s 4618 16200 4674 17000 0 FreeSans 224 90 0 0 gpio_defaults[8]
port 11 nsew signal input
flabel metal2 s 5078 16200 5134 17000 0 FreeSans 224 90 0 0 gpio_defaults[9]
port 12 nsew signal input
flabel metal3 s 14000 4824 34000 4944 0 FreeSans 480 0 0 0 mgmt_gpio_in
port 13 nsew signal tristate
flabel metal3 s 14000 5640 34000 5760 0 FreeSans 480 0 0 0 mgmt_gpio_oeb
port 14 nsew signal input
flabel metal3 s 14000 6048 34000 6168 0 FreeSans 480 0 0 0 mgmt_gpio_out
port 15 nsew signal input
flabel metal3 s 14000 5232 34000 5352 0 FreeSans 480 0 0 0 one
port 16 nsew signal tristate
flabel metal3 s 14000 6456 34000 6576 0 FreeSans 480 0 0 0 pad_gpio_ana_en
port 17 nsew signal tristate
flabel metal3 s 14000 6864 34000 6984 0 FreeSans 480 0 0 0 pad_gpio_ana_pol
port 18 nsew signal tristate
flabel metal3 s 14000 7272 34000 7392 0 FreeSans 480 0 0 0 pad_gpio_ana_sel
port 19 nsew signal tristate
flabel metal3 s 14000 7680 34000 7800 0 FreeSans 480 0 0 0 pad_gpio_dm[0]
port 20 nsew signal tristate
flabel metal3 s 14000 8088 34000 8208 0 FreeSans 480 0 0 0 pad_gpio_dm[1]
port 21 nsew signal tristate
flabel metal3 s 14000 8496 34000 8616 0 FreeSans 480 0 0 0 pad_gpio_dm[2]
port 22 nsew signal tristate
flabel metal3 s 14000 8904 34000 9024 0 FreeSans 480 0 0 0 pad_gpio_holdover
port 23 nsew signal tristate
flabel metal3 s 14000 9312 34000 9432 0 FreeSans 480 0 0 0 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
flabel metal3 s 14000 9720 34000 9840 0 FreeSans 480 0 0 0 pad_gpio_in
port 25 nsew signal input
flabel metal3 s 14000 10128 34000 10248 0 FreeSans 480 0 0 0 pad_gpio_inenb
port 26 nsew signal tristate
flabel metal3 s 14000 10536 34000 10656 0 FreeSans 480 0 0 0 pad_gpio_out
port 27 nsew signal tristate
flabel metal3 s 14000 10944 34000 11064 0 FreeSans 480 0 0 0 pad_gpio_outenb
port 28 nsew signal tristate
flabel metal3 s 14000 11352 34000 11472 0 FreeSans 480 0 0 0 pad_gpio_slow_sel
port 29 nsew signal tristate
flabel metal3 s 14000 11760 34000 11880 0 FreeSans 480 0 0 0 pad_gpio_vtrip_sel
port 30 nsew signal tristate
flabel metal3 s 14000 12168 34000 12288 0 FreeSans 480 0 0 0 resetn
port 31 nsew signal input
flabel metal3 s 14000 12576 34000 12696 0 FreeSans 480 0 0 0 resetn_out
port 32 nsew signal tristate
flabel metal3 s 14000 12984 34000 13104 0 FreeSans 480 0 0 0 serial_clock
port 33 nsew signal input
flabel metal3 s 14000 13392 34000 13512 0 FreeSans 480 0 0 0 serial_clock_out
port 34 nsew signal tristate
flabel metal3 s 14000 13800 34000 13920 0 FreeSans 480 0 0 0 serial_data_in
port 35 nsew signal input
flabel metal3 s 14000 14208 34000 14328 0 FreeSans 480 0 0 0 serial_data_out
port 36 nsew signal tristate
flabel metal3 s 14000 14616 34000 14736 0 FreeSans 480 0 0 0 serial_load
port 37 nsew signal input
flabel metal3 s 14000 15024 34000 15144 0 FreeSans 480 0 0 0 serial_load_out
port 38 nsew signal tristate
flabel metal3 s 14000 15432 34000 15552 0 FreeSans 480 0 0 0 user_gpio_in
port 39 nsew signal tristate
flabel metal3 s 14000 15840 34000 15960 0 FreeSans 480 0 0 0 user_gpio_oeb
port 40 nsew signal input
flabel metal3 s 14000 16248 34000 16368 0 FreeSans 480 0 0 0 user_gpio_out
port 41 nsew signal input
flabel metal4 s 2560 4893 2880 15824 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 7560 928 7880 15824 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 928 9892 1248 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 4928 9892 5248 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 8928 9892 9248 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 12928 9892 13248 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 4560 1040 4880 15824 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 2928 9892 3248 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 3560 1040 3880 15824 0 FreeSans 1920 90 0 0 vssd
port 44 nsew ground bidirectional
flabel metal4 s 8560 1040 8880 15824 0 FreeSans 1920 90 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 1928 9892 2248 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 5928 9892 6248 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 9928 9892 10248 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 13928 9892 14248 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal4 s 5560 1040 5880 15824 0 FreeSans 1920 90 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 3928 9892 4248 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal3 s 14000 4416 34000 4536 0 FreeSans 480 0 0 0 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 17000
<< end >>
