magic
tech sky130A
magscale 1 2
timestamp 1664316539
<< obsli1 >>
rect 0 0 33962 17000
<< obsm1 >>
rect 106 0 34000 17000
<< metal2 >>
rect 938 16200 994 17000
rect 1398 16200 1454 17000
rect 1858 16200 1914 17000
rect 2318 16200 2374 17000
rect 2778 16200 2834 17000
rect 3238 16200 3294 17000
rect 3698 16200 3754 17000
rect 4158 16200 4214 17000
rect 4618 16200 4674 17000
rect 5078 16200 5134 17000
rect 5538 16200 5594 17000
rect 5998 16200 6054 17000
rect 6458 16200 6514 17000
<< obsm2 >>
rect 112 16144 882 17000
rect 1050 16144 1342 17000
rect 1510 16144 1802 17000
rect 1970 16144 2262 17000
rect 2430 16144 2722 17000
rect 2890 16144 3182 17000
rect 3350 16144 3642 17000
rect 3810 16144 4102 17000
rect 4270 16144 4562 17000
rect 4730 16144 5022 17000
rect 5190 16144 5482 17000
rect 5650 16144 5942 17000
rect 6110 16144 6402 17000
rect 6570 16144 34000 17000
rect 112 0 34000 16144
<< metal3 >>
rect 14000 16248 34000 16368
rect 14000 15840 34000 15960
rect 14000 15432 34000 15552
rect 14000 15024 34000 15144
rect 14000 14616 34000 14736
rect 14000 14208 34000 14328
rect 14000 13800 34000 13920
rect 14000 13392 34000 13512
rect 14000 12984 34000 13104
rect 14000 12576 34000 12696
rect 14000 12168 34000 12288
rect 14000 11760 34000 11880
rect 14000 11352 34000 11472
rect 14000 10944 34000 11064
rect 14000 10536 34000 10656
rect 14000 10128 34000 10248
rect 14000 9720 34000 9840
rect 14000 9312 34000 9432
rect 14000 8904 34000 9024
rect 14000 8496 34000 8616
rect 14000 8088 34000 8208
rect 14000 7680 34000 7800
rect 14000 7272 34000 7392
rect 14000 6864 34000 6984
rect 14000 6456 34000 6576
rect 14000 6048 34000 6168
rect 14000 5640 34000 5760
rect 14000 5232 34000 5352
rect 14000 4824 34000 4944
rect 14000 4416 34000 4536
<< obsm3 >>
rect 197 16448 16866 16557
rect 197 16168 13920 16448
rect 197 16040 16866 16168
rect 197 15760 13920 16040
rect 197 15632 16866 15760
rect 197 15352 13920 15632
rect 197 15224 16866 15352
rect 197 14944 13920 15224
rect 197 14816 16866 14944
rect 197 14536 13920 14816
rect 197 14408 16866 14536
rect 197 14128 13920 14408
rect 197 14000 16866 14128
rect 197 13720 13920 14000
rect 197 13592 16866 13720
rect 197 13312 13920 13592
rect 197 13184 16866 13312
rect 197 12904 13920 13184
rect 197 12776 16866 12904
rect 197 12496 13920 12776
rect 197 12368 16866 12496
rect 197 12088 13920 12368
rect 197 11960 16866 12088
rect 197 11680 13920 11960
rect 197 11552 16866 11680
rect 197 11272 13920 11552
rect 197 11144 16866 11272
rect 197 10864 13920 11144
rect 197 10736 16866 10864
rect 197 10456 13920 10736
rect 197 10328 16866 10456
rect 197 10048 13920 10328
rect 197 9920 16866 10048
rect 197 9640 13920 9920
rect 197 9512 16866 9640
rect 197 9232 13920 9512
rect 197 9104 16866 9232
rect 197 8824 13920 9104
rect 197 8696 16866 8824
rect 197 8416 13920 8696
rect 197 8288 16866 8416
rect 197 8008 13920 8288
rect 197 7880 16866 8008
rect 197 7600 13920 7880
rect 197 7472 16866 7600
rect 197 7192 13920 7472
rect 197 7064 16866 7192
rect 197 6784 13920 7064
rect 197 6656 16866 6784
rect 197 6376 13920 6656
rect 197 6248 16866 6376
rect 197 5968 13920 6248
rect 197 5840 16866 5968
rect 197 5560 13920 5840
rect 197 5432 16866 5560
rect 197 5152 13920 5432
rect 197 5024 16866 5152
rect 197 4744 13920 5024
rect 197 4616 16866 4744
rect 197 4336 13920 4616
rect 197 35 16866 4336
<< metal4 >>
rect 2560 4893 2880 15824
rect 3560 1040 3880 15824
rect 4560 1040 4880 15824
rect 5560 1040 5880 15824
rect 7560 928 7880 15824
rect 8560 1040 8880 15824
<< obsm4 >>
rect 0 15904 34000 17000
rect 0 4813 2480 15904
rect 2960 4813 3480 15904
rect 0 960 3480 4813
rect 3960 960 4480 15904
rect 4960 960 5480 15904
rect 5960 960 7480 15904
rect 0 848 7480 960
rect 7960 960 8480 15904
rect 8960 960 34000 15904
rect 7960 848 34000 960
rect 0 0 34000 848
<< metal5 >>
rect 872 13928 9892 14248
rect 872 12928 9892 13248
rect 872 9928 9892 10248
rect 872 8928 9892 9248
rect 872 5928 9892 6248
rect 872 4928 9892 5248
rect 872 3928 9892 4248
rect 872 2928 9892 3248
rect 872 1928 9892 2248
rect 872 928 9892 1248
<< obsm5 >>
rect 2140 14568 34000 17000
rect 10212 13608 34000 14568
rect 2140 13568 34000 13608
rect 10212 12608 34000 13568
rect 2140 10568 34000 12608
rect 10212 9608 34000 10568
rect 2140 9568 34000 9608
rect 10212 8608 34000 9568
rect 2140 6568 34000 8608
rect 10212 5608 34000 6568
rect 2140 5568 34000 5608
rect 10212 4608 34000 5568
rect 2140 4568 34000 4608
rect 10212 3608 34000 4568
rect 2140 3568 34000 3608
rect 10212 2608 34000 3568
rect 2140 2568 34000 2608
rect 10212 1608 34000 2568
rect 2140 1568 34000 1608
rect 10212 608 34000 1568
rect 2140 0 34000 608
<< labels >>
rlabel metal2 s 938 16200 994 17000 6 gpio_defaults[0]
port 1 nsew signal input
rlabel metal2 s 5538 16200 5594 17000 6 gpio_defaults[10]
port 2 nsew signal input
rlabel metal2 s 5998 16200 6054 17000 6 gpio_defaults[11]
port 3 nsew signal input
rlabel metal2 s 6458 16200 6514 17000 6 gpio_defaults[12]
port 4 nsew signal input
rlabel metal2 s 1398 16200 1454 17000 6 gpio_defaults[1]
port 5 nsew signal input
rlabel metal2 s 1858 16200 1914 17000 6 gpio_defaults[2]
port 6 nsew signal input
rlabel metal2 s 2318 16200 2374 17000 6 gpio_defaults[3]
port 7 nsew signal input
rlabel metal2 s 2778 16200 2834 17000 6 gpio_defaults[4]
port 8 nsew signal input
rlabel metal2 s 3238 16200 3294 17000 6 gpio_defaults[5]
port 9 nsew signal input
rlabel metal2 s 3698 16200 3754 17000 6 gpio_defaults[6]
port 10 nsew signal input
rlabel metal2 s 4158 16200 4214 17000 6 gpio_defaults[7]
port 11 nsew signal input
rlabel metal2 s 4618 16200 4674 17000 6 gpio_defaults[8]
port 12 nsew signal input
rlabel metal2 s 5078 16200 5134 17000 6 gpio_defaults[9]
port 13 nsew signal input
rlabel metal3 s 14000 4824 34000 4944 6 mgmt_gpio_in
port 14 nsew signal output
rlabel metal3 s 14000 5640 34000 5760 6 mgmt_gpio_oeb
port 15 nsew signal input
rlabel metal3 s 14000 6048 34000 6168 6 mgmt_gpio_out
port 16 nsew signal input
rlabel metal3 s 14000 5232 34000 5352 6 one
port 17 nsew signal output
rlabel metal3 s 14000 6456 34000 6576 6 pad_gpio_ana_en
port 18 nsew signal output
rlabel metal3 s 14000 6864 34000 6984 6 pad_gpio_ana_pol
port 19 nsew signal output
rlabel metal3 s 14000 7272 34000 7392 6 pad_gpio_ana_sel
port 20 nsew signal output
rlabel metal3 s 14000 7680 34000 7800 6 pad_gpio_dm[0]
port 21 nsew signal output
rlabel metal3 s 14000 8088 34000 8208 6 pad_gpio_dm[1]
port 22 nsew signal output
rlabel metal3 s 14000 8496 34000 8616 6 pad_gpio_dm[2]
port 23 nsew signal output
rlabel metal3 s 14000 8904 34000 9024 6 pad_gpio_holdover
port 24 nsew signal output
rlabel metal3 s 14000 9312 34000 9432 6 pad_gpio_ib_mode_sel
port 25 nsew signal output
rlabel metal3 s 14000 9720 34000 9840 6 pad_gpio_in
port 26 nsew signal input
rlabel metal3 s 14000 10128 34000 10248 6 pad_gpio_inenb
port 27 nsew signal output
rlabel metal3 s 14000 10536 34000 10656 6 pad_gpio_out
port 28 nsew signal output
rlabel metal3 s 14000 10944 34000 11064 6 pad_gpio_outenb
port 29 nsew signal output
rlabel metal3 s 14000 11352 34000 11472 6 pad_gpio_slow_sel
port 30 nsew signal output
rlabel metal3 s 14000 11760 34000 11880 6 pad_gpio_vtrip_sel
port 31 nsew signal output
rlabel metal3 s 14000 12168 34000 12288 6 resetn
port 32 nsew signal input
rlabel metal3 s 14000 12576 34000 12696 6 resetn_out
port 33 nsew signal output
rlabel metal3 s 14000 12984 34000 13104 6 serial_clock
port 34 nsew signal input
rlabel metal3 s 14000 13392 34000 13512 6 serial_clock_out
port 35 nsew signal output
rlabel metal3 s 14000 13800 34000 13920 6 serial_data_in
port 36 nsew signal input
rlabel metal3 s 14000 14208 34000 14328 6 serial_data_out
port 37 nsew signal output
rlabel metal3 s 14000 14616 34000 14736 6 serial_load
port 38 nsew signal input
rlabel metal3 s 14000 15024 34000 15144 6 serial_load_out
port 39 nsew signal output
rlabel metal3 s 14000 15432 34000 15552 6 user_gpio_in
port 40 nsew signal output
rlabel metal3 s 14000 15840 34000 15960 6 user_gpio_oeb
port 41 nsew signal input
rlabel metal3 s 14000 16248 34000 16368 6 user_gpio_out
port 42 nsew signal input
rlabel metal4 s 2560 4893 2880 15824 6 vccd
port 43 nsew power bidirectional
rlabel metal4 s 7560 928 7880 15824 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 928 9892 1248 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 4928 9892 5248 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 8928 9892 9248 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 12928 9892 13248 6 vccd
port 43 nsew power bidirectional
rlabel metal4 s 4560 1040 4880 15824 6 vccd1
port 44 nsew power bidirectional
rlabel metal5 s 872 2928 9892 3248 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 3560 1040 3880 15824 6 vssd
port 45 nsew ground bidirectional
rlabel metal4 s 8560 1040 8880 15824 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s 872 1928 9892 2248 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s 872 5928 9892 6248 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s 872 9928 9892 10248 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s 872 13928 9892 14248 6 vssd
port 45 nsew ground bidirectional
rlabel metal4 s 5560 1040 5880 15824 6 vssd1
port 46 nsew ground bidirectional
rlabel metal5 s 872 3928 9892 4248 6 vssd1
port 46 nsew ground bidirectional
rlabel metal3 s 14000 4416 34000 4536 6 zero
port 47 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 34000 17000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 706176
string GDS_FILE /openlane/designs/gpio_control_block/runs/RUN_6/results/signoff/gpio_control_block.magic.gds
string GDS_START 185666
<< end >>

