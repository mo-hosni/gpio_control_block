magic
tech sky130A
magscale 1 2
timestamp 1664190901
<< obsli1 >>
rect 0 0 33962 17000
<< obsm1 >>
rect 106 0 34000 17000
<< metal2 >>
rect 938 16200 994 17000
rect 1398 16200 1454 17000
rect 1858 16200 1914 17000
rect 2318 16200 2374 17000
rect 2778 16200 2834 17000
rect 3238 16200 3294 17000
rect 3698 16200 3754 17000
rect 4158 16200 4214 17000
rect 4618 16200 4674 17000
rect 5078 16200 5134 17000
rect 5538 16200 5594 17000
rect 5998 16200 6054 17000
rect 6458 16200 6514 17000
<< obsm2 >>
rect 18 16144 882 17000
rect 1050 16144 1342 17000
rect 1510 16144 1802 17000
rect 1970 16144 2262 17000
rect 2430 16144 2722 17000
rect 2890 16144 3182 17000
rect 3350 16144 3642 17000
rect 3810 16144 4102 17000
rect 4270 16144 4562 17000
rect 4730 16144 5022 17000
rect 5190 16144 5482 17000
rect 5650 16144 5942 17000
rect 6110 16144 6402 17000
rect 6570 16144 34000 17000
rect 18 0 34000 16144
<< metal3 >>
rect 14000 16328 34000 16448
rect 14000 15920 34000 16040
rect 14000 15512 34000 15632
rect 14000 15104 34000 15224
rect 14000 14696 34000 14816
rect 14000 14288 34000 14408
rect 14000 13880 34000 14000
rect 14000 13472 34000 13592
rect 14000 13064 34000 13184
rect 14000 12656 34000 12776
rect 14000 12248 34000 12368
rect 14000 11840 34000 11960
rect 14000 11432 34000 11552
rect 14000 11024 34000 11144
rect 14000 10616 34000 10736
rect 14000 10208 34000 10328
rect 14000 9800 34000 9920
rect 14000 9392 34000 9512
rect 14000 8984 34000 9104
rect 14000 8576 34000 8696
rect 14000 8168 34000 8288
rect 14000 7760 34000 7880
rect 14000 7352 34000 7472
rect 14000 6944 34000 7064
rect 14000 6536 34000 6656
rect 14000 6128 34000 6248
rect 14000 5720 34000 5840
rect 14000 5312 34000 5432
rect 14000 4904 34000 5024
rect 14000 4496 34000 4616
<< obsm3 >>
rect 13 16528 17099 16965
rect 13 16248 13920 16528
rect 13 16120 17099 16248
rect 13 15840 13920 16120
rect 13 15712 17099 15840
rect 13 15432 13920 15712
rect 13 15304 17099 15432
rect 13 15024 13920 15304
rect 13 14896 17099 15024
rect 13 14616 13920 14896
rect 13 14488 17099 14616
rect 13 14208 13920 14488
rect 13 14080 17099 14208
rect 13 13800 13920 14080
rect 13 13672 17099 13800
rect 13 13392 13920 13672
rect 13 13264 17099 13392
rect 13 12984 13920 13264
rect 13 12856 17099 12984
rect 13 12576 13920 12856
rect 13 12448 17099 12576
rect 13 12168 13920 12448
rect 13 12040 17099 12168
rect 13 11760 13920 12040
rect 13 11632 17099 11760
rect 13 11352 13920 11632
rect 13 11224 17099 11352
rect 13 10944 13920 11224
rect 13 10816 17099 10944
rect 13 10536 13920 10816
rect 13 10408 17099 10536
rect 13 10128 13920 10408
rect 13 10000 17099 10128
rect 13 9720 13920 10000
rect 13 9592 17099 9720
rect 13 9312 13920 9592
rect 13 9184 17099 9312
rect 13 8904 13920 9184
rect 13 8776 17099 8904
rect 13 8496 13920 8776
rect 13 8368 17099 8496
rect 13 8088 13920 8368
rect 13 7960 17099 8088
rect 13 7680 13920 7960
rect 13 7552 17099 7680
rect 13 7272 13920 7552
rect 13 7144 17099 7272
rect 13 6864 13920 7144
rect 13 6736 17099 6864
rect 13 6456 13920 6736
rect 13 6328 17099 6456
rect 13 6048 13920 6328
rect 13 5920 17099 6048
rect 13 5640 13920 5920
rect 13 5512 17099 5640
rect 13 5232 13920 5512
rect 13 5104 17099 5232
rect 13 4824 13920 5104
rect 13 4696 17099 4824
rect 13 4416 13920 4696
rect 13 171 17099 4416
<< metal4 >>
rect 2560 4893 2880 15824
rect 3560 1040 3880 15824
rect 4560 1040 4880 15824
rect 5560 1040 5880 15824
rect 7560 928 7880 15824
rect 8560 1040 8880 15824
rect 9560 1040 9880 15824
<< obsm4 >>
rect 59 15904 34000 17000
rect 59 4813 2480 15904
rect 2960 4813 3480 15904
rect 59 960 3480 4813
rect 3960 960 4480 15904
rect 4960 960 5480 15904
rect 5960 960 7480 15904
rect 59 848 7480 960
rect 7960 960 8480 15904
rect 8960 960 9480 15904
rect 9960 960 34000 15904
rect 7960 848 34000 960
rect 59 0 34000 848
<< metal5 >>
rect 872 14928 9892 15248
rect 872 13928 9892 14248
rect 872 12928 9892 13248
rect 872 10928 9892 11248
rect 872 9928 9892 10248
rect 872 8928 9892 9248
rect 872 6928 9892 7248
rect 872 5928 9892 6248
rect 872 4928 9892 5248
rect 872 3928 9892 4248
rect 872 2928 9892 3248
rect 872 1928 9892 2248
rect 872 928 9892 1248
<< obsm5 >>
rect 13400 0 34000 17000
<< labels >>
rlabel metal2 s 938 16200 994 17000 6 gpio_defaults[0]
port 1 nsew signal input
rlabel metal2 s 5538 16200 5594 17000 6 gpio_defaults[10]
port 2 nsew signal input
rlabel metal2 s 5998 16200 6054 17000 6 gpio_defaults[11]
port 3 nsew signal input
rlabel metal2 s 6458 16200 6514 17000 6 gpio_defaults[12]
port 4 nsew signal input
rlabel metal2 s 1398 16200 1454 17000 6 gpio_defaults[1]
port 5 nsew signal input
rlabel metal2 s 1858 16200 1914 17000 6 gpio_defaults[2]
port 6 nsew signal input
rlabel metal2 s 2318 16200 2374 17000 6 gpio_defaults[3]
port 7 nsew signal input
rlabel metal2 s 2778 16200 2834 17000 6 gpio_defaults[4]
port 8 nsew signal input
rlabel metal2 s 3238 16200 3294 17000 6 gpio_defaults[5]
port 9 nsew signal input
rlabel metal2 s 3698 16200 3754 17000 6 gpio_defaults[6]
port 10 nsew signal input
rlabel metal2 s 4158 16200 4214 17000 6 gpio_defaults[7]
port 11 nsew signal input
rlabel metal2 s 4618 16200 4674 17000 6 gpio_defaults[8]
port 12 nsew signal input
rlabel metal2 s 5078 16200 5134 17000 6 gpio_defaults[9]
port 13 nsew signal input
rlabel metal3 s 14000 4904 34000 5024 6 mgmt_gpio_in
port 14 nsew signal output
rlabel metal3 s 14000 5720 34000 5840 6 mgmt_gpio_oeb
port 15 nsew signal input
rlabel metal3 s 14000 6128 34000 6248 6 mgmt_gpio_out
port 16 nsew signal input
rlabel metal3 s 14000 5312 34000 5432 6 one
port 17 nsew signal output
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_ana_en
port 18 nsew signal output
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_ana_pol
port 19 nsew signal output
rlabel metal3 s 14000 7352 34000 7472 6 pad_gpio_ana_sel
port 20 nsew signal output
rlabel metal3 s 14000 7760 34000 7880 6 pad_gpio_dm[0]
port 21 nsew signal output
rlabel metal3 s 14000 8168 34000 8288 6 pad_gpio_dm[1]
port 22 nsew signal output
rlabel metal3 s 14000 8576 34000 8696 6 pad_gpio_dm[2]
port 23 nsew signal output
rlabel metal3 s 14000 8984 34000 9104 6 pad_gpio_holdover
port 24 nsew signal output
rlabel metal3 s 14000 9392 34000 9512 6 pad_gpio_ib_mode_sel
port 25 nsew signal output
rlabel metal3 s 14000 9800 34000 9920 6 pad_gpio_in
port 26 nsew signal input
rlabel metal3 s 14000 10208 34000 10328 6 pad_gpio_inenb
port 27 nsew signal output
rlabel metal3 s 14000 10616 34000 10736 6 pad_gpio_out
port 28 nsew signal output
rlabel metal3 s 14000 11024 34000 11144 6 pad_gpio_outenb
port 29 nsew signal output
rlabel metal3 s 14000 11432 34000 11552 6 pad_gpio_slow_sel
port 30 nsew signal output
rlabel metal3 s 14000 11840 34000 11960 6 pad_gpio_vtrip_sel
port 31 nsew signal output
rlabel metal3 s 14000 12248 34000 12368 6 resetn
port 32 nsew signal input
rlabel metal3 s 14000 12656 34000 12776 6 resetn_out
port 33 nsew signal output
rlabel metal3 s 14000 13064 34000 13184 6 serial_clock
port 34 nsew signal input
rlabel metal3 s 14000 13472 34000 13592 6 serial_clock_out
port 35 nsew signal output
rlabel metal3 s 14000 13880 34000 14000 6 serial_data_in
port 36 nsew signal input
rlabel metal3 s 14000 14288 34000 14408 6 serial_data_out
port 37 nsew signal output
rlabel metal3 s 14000 14696 34000 14816 6 serial_load
port 38 nsew signal input
rlabel metal3 s 14000 15104 34000 15224 6 serial_load_out
port 39 nsew signal output
rlabel metal3 s 14000 15512 34000 15632 6 user_gpio_in
port 40 nsew signal output
rlabel metal3 s 14000 15920 34000 16040 6 user_gpio_oeb
port 41 nsew signal input
rlabel metal3 s 14000 16328 34000 16448 6 user_gpio_out
port 42 nsew signal input
rlabel metal4 s 2560 4893 2880 15824 6 vccd
port 43 nsew power bidirectional
rlabel metal4 s 7560 928 7880 15824 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 928 9892 1248 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 4928 9892 5248 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 8928 9892 9248 6 vccd
port 43 nsew power bidirectional
rlabel metal5 s 872 12928 9892 13248 6 vccd
port 43 nsew power bidirectional
rlabel metal4 s 4560 1040 4880 15824 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 9560 1040 9880 15824 6 vccd1
port 44 nsew power bidirectional
rlabel metal5 s 872 2928 9892 3248 6 vccd1
port 44 nsew power bidirectional
rlabel metal5 s 872 6928 9892 7248 6 vccd1
port 44 nsew power bidirectional
rlabel metal5 s 872 10928 9892 11248 6 vccd1
port 44 nsew power bidirectional
rlabel metal5 s 872 14928 9892 15248 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 3560 1040 3880 15824 6 vssd
port 45 nsew ground bidirectional
rlabel metal4 s 8560 1040 8880 15824 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s 872 1928 9892 2248 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s 872 5928 9892 6248 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s 872 9928 9892 10248 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s 872 13928 9892 14248 6 vssd
port 45 nsew ground bidirectional
rlabel metal4 s 5560 1040 5880 15824 6 vssd1
port 46 nsew ground bidirectional
rlabel metal5 s 872 3928 9892 4248 6 vssd1
port 46 nsew ground bidirectional
rlabel metal3 s 14000 4496 34000 4616 6 zero
port 47 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 34000 17000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 686962
string GDS_FILE /openlane/designs/gpio_control_block/runs/RUN_27/results/signoff/gpio_control_block.magic.gds
string GDS_START 185666
<< end >>

