magic
tech sky130A
magscale 1 2
timestamp 1664190920
<< checkpaint >>
rect -3919 -3765 37932 20932
<< viali >>
rect 2329 15657 2363 15691
rect 5733 15657 5767 15691
rect 4721 15521 4755 15555
rect 1777 15453 1811 15487
rect 2513 15453 2547 15487
rect 3249 15453 3283 15487
rect 4997 15453 5031 15487
rect 5549 15453 5583 15487
rect 8401 15453 8435 15487
rect 8953 15453 8987 15487
rect 2973 15385 3007 15419
rect 3157 15385 3191 15419
rect 8125 15385 8159 15419
rect 1593 15317 1627 15351
rect 3065 15317 3099 15351
rect 6653 15317 6687 15351
rect 9137 15317 9171 15351
rect 6653 15113 6687 15147
rect 1501 15045 1535 15079
rect 2605 15045 2639 15079
rect 3433 15045 3467 15079
rect 8125 15045 8159 15079
rect 1685 14977 1719 15011
rect 2421 14977 2455 15011
rect 3249 14977 3283 15011
rect 4077 14977 4111 15011
rect 5733 14977 5767 15011
rect 8953 14977 8987 15011
rect 8401 14909 8435 14943
rect 2789 14841 2823 14875
rect 5181 14841 5215 14875
rect 1869 14773 1903 14807
rect 3617 14773 3651 14807
rect 4721 14773 4755 14807
rect 9137 14773 9171 14807
rect 2973 14433 3007 14467
rect 4813 14433 4847 14467
rect 5273 14433 5307 14467
rect 3249 14365 3283 14399
rect 3985 14365 4019 14399
rect 7757 14365 7791 14399
rect 8953 14365 8987 14399
rect 4445 14297 4479 14331
rect 4629 14297 4663 14331
rect 7021 14297 7055 14331
rect 9137 14297 9171 14331
rect 1501 14229 1535 14263
rect 3893 14229 3927 14263
rect 8309 14229 8343 14263
rect 9321 14229 9355 14263
rect 2605 14025 2639 14059
rect 5457 14025 5491 14059
rect 6653 14025 6687 14059
rect 1593 13889 1627 13923
rect 3065 13889 3099 13923
rect 4537 13889 4571 13923
rect 5641 13889 5675 13923
rect 5825 13889 5859 13923
rect 7113 13889 7147 13923
rect 8585 13889 8619 13923
rect 8953 13889 8987 13923
rect 2145 13821 2179 13855
rect 4905 13821 4939 13855
rect 4445 13345 4479 13379
rect 7481 13345 7515 13379
rect 3893 13277 3927 13311
rect 5181 13277 5215 13311
rect 5549 13277 5583 13311
rect 7021 13277 7055 13311
rect 8033 13277 8067 13311
rect 8953 13277 8987 13311
rect 1501 13209 1535 13243
rect 2789 13141 2823 13175
rect 8217 13141 8251 13175
rect 9137 13141 9171 13175
rect 8309 12937 8343 12971
rect 1593 12801 1627 12835
rect 2973 12801 3007 12835
rect 4445 12801 4479 12835
rect 5365 12801 5399 12835
rect 6561 12801 6595 12835
rect 9229 12801 9263 12835
rect 2605 12733 2639 12767
rect 5641 12733 5675 12767
rect 6837 12733 6871 12767
rect 2145 12597 2179 12631
rect 4905 12597 4939 12631
rect 9137 12597 9171 12631
rect 2973 12257 3007 12291
rect 7481 12257 7515 12291
rect 3249 12189 3283 12223
rect 3801 12189 3835 12223
rect 3985 12189 4019 12223
rect 4445 12189 4479 12223
rect 4813 12189 4847 12223
rect 6285 12189 6319 12223
rect 8953 12189 8987 12223
rect 9137 12121 9171 12155
rect 1501 12053 1535 12087
rect 3893 12053 3927 12087
rect 6745 12053 6779 12087
rect 8125 12053 8159 12087
rect 9321 12053 9355 12087
rect 8125 11849 8159 11883
rect 9229 11849 9263 11883
rect 5825 11781 5859 11815
rect 8861 11781 8895 11815
rect 3617 11713 3651 11747
rect 6377 11713 6411 11747
rect 8769 11713 8803 11747
rect 9045 11713 9079 11747
rect 3341 11645 3375 11679
rect 4169 11645 4203 11679
rect 6653 11645 6687 11679
rect 1869 11509 1903 11543
rect 3249 11305 3283 11339
rect 1593 11169 1627 11203
rect 2605 11169 2639 11203
rect 4905 11169 4939 11203
rect 8033 11169 8067 11203
rect 7665 11101 7699 11135
rect 8953 11101 8987 11135
rect 2145 11033 2179 11067
rect 4261 11033 4295 11067
rect 5549 11033 5583 11067
rect 7205 11033 7239 11067
rect 7849 11033 7883 11067
rect 9137 10965 9171 10999
rect 4813 10761 4847 10795
rect 1409 10693 1443 10727
rect 5457 10693 5491 10727
rect 1593 10625 1627 10659
rect 2881 10625 2915 10659
rect 4353 10625 4387 10659
rect 5641 10625 5675 10659
rect 6837 10625 6871 10659
rect 8309 10625 8343 10659
rect 9137 10625 9171 10659
rect 2513 10557 2547 10591
rect 8677 10557 8711 10591
rect 9229 10557 9263 10591
rect 1777 10421 1811 10455
rect 5825 10421 5859 10455
rect 6377 10421 6411 10455
rect 2145 10217 2179 10251
rect 8953 10217 8987 10251
rect 9137 10217 9171 10251
rect 1593 10081 1627 10115
rect 2605 10081 2639 10115
rect 4077 10081 4111 10115
rect 8309 10081 8343 10115
rect 3801 10013 3835 10047
rect 6009 10013 6043 10047
rect 6377 10013 6411 10047
rect 7849 10013 7883 10047
rect 9321 9945 9355 9979
rect 3249 9877 3283 9911
rect 5549 9877 5583 9911
rect 8033 9877 8067 9911
rect 9121 9877 9155 9911
rect 7389 9605 7423 9639
rect 9137 9605 9171 9639
rect 3065 9537 3099 9571
rect 3525 9537 3559 9571
rect 5365 9537 5399 9571
rect 6469 9537 6503 9571
rect 1501 9469 1535 9503
rect 2697 9469 2731 9503
rect 3893 9469 3927 9503
rect 5825 9469 5859 9503
rect 6561 9333 6595 9367
rect 6929 9333 6963 9367
rect 4721 9129 4755 9163
rect 1777 8993 1811 9027
rect 4077 8993 4111 9027
rect 7665 8993 7699 9027
rect 1501 8925 1535 8959
rect 5273 8925 5307 8959
rect 7481 8925 7515 8959
rect 9045 8925 9079 8959
rect 3249 8789 3283 8823
rect 6561 8789 6595 8823
rect 9137 8789 9171 8823
rect 5089 8585 5123 8619
rect 5641 8585 5675 8619
rect 6377 8585 6411 8619
rect 9137 8517 9171 8551
rect 1777 8449 1811 8483
rect 2329 8449 2363 8483
rect 3157 8449 3191 8483
rect 4629 8449 4663 8483
rect 5825 8449 5859 8483
rect 6929 8449 6963 8483
rect 9321 8449 9355 8483
rect 2789 8381 2823 8415
rect 8217 8381 8251 8415
rect 3801 7905 3835 7939
rect 1501 7837 1535 7871
rect 7021 7837 7055 7871
rect 8033 7837 8067 7871
rect 9137 7837 9171 7871
rect 3249 7769 3283 7803
rect 5273 7769 5307 7803
rect 8953 7769 8987 7803
rect 4445 7701 4479 7735
rect 7481 7701 7515 7735
rect 9321 7701 9355 7735
rect 5825 7497 5859 7531
rect 9137 7497 9171 7531
rect 1869 7429 1903 7463
rect 3617 7429 3651 7463
rect 4353 7429 4387 7463
rect 8217 7361 8251 7395
rect 9321 7361 9355 7395
rect 4077 7293 4111 7327
rect 6377 7293 6411 7327
rect 6745 7293 6779 7327
rect 8677 7157 8711 7191
rect 1501 6817 1535 6851
rect 1777 6817 1811 6851
rect 3893 6817 3927 6851
rect 5641 6749 5675 6783
rect 6101 6749 6135 6783
rect 6469 6749 6503 6783
rect 7941 6749 7975 6783
rect 8953 6749 8987 6783
rect 5365 6681 5399 6715
rect 9137 6681 9171 6715
rect 3249 6613 3283 6647
rect 8401 6613 8435 6647
rect 9321 6613 9355 6647
rect 2329 6409 2363 6443
rect 3249 6409 3283 6443
rect 4997 6273 5031 6307
rect 5825 6273 5859 6307
rect 6929 6273 6963 6307
rect 8401 6273 8435 6307
rect 1777 6205 1811 6239
rect 4721 6205 4755 6239
rect 6561 6205 6595 6239
rect 5641 6137 5675 6171
rect 8861 6069 8895 6103
rect 2513 5865 2547 5899
rect 5549 5865 5583 5899
rect 7021 5865 7055 5899
rect 8309 5865 8343 5899
rect 1777 5797 1811 5831
rect 3801 5729 3835 5763
rect 6377 5729 6411 5763
rect 1961 5661 1995 5695
rect 2697 5661 2731 5695
rect 7757 5661 7791 5695
rect 8401 5661 8435 5695
rect 9229 5661 9263 5695
rect 4077 5593 4111 5627
rect 8953 5593 8987 5627
rect 9137 5593 9171 5627
rect 7573 5525 7607 5559
rect 9045 5525 9079 5559
rect 4077 5321 4111 5355
rect 5825 5321 5859 5355
rect 7297 5321 7331 5355
rect 9229 5253 9263 5287
rect 4169 5185 4203 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 7205 5185 7239 5219
rect 9137 5185 9171 5219
rect 5181 5117 5215 5151
rect 6745 4981 6779 5015
rect 3617 4777 3651 4811
rect 4721 4777 4755 4811
rect 5273 4777 5307 4811
rect 6745 4777 6779 4811
rect 7389 4777 7423 4811
rect 8401 4777 8435 4811
rect 9229 4777 9263 4811
rect 6009 4709 6043 4743
rect 3525 4573 3559 4607
rect 4537 4573 4571 4607
rect 5181 4573 5215 4607
rect 5365 4573 5399 4607
rect 6193 4573 6227 4607
rect 6837 4573 6871 4607
rect 7297 4573 7331 4607
rect 7481 4573 7515 4607
rect 8585 4573 8619 4607
rect 9045 4573 9079 4607
rect 7021 4233 7055 4267
rect 7573 4233 7607 4267
rect 3709 4097 3743 4131
rect 4077 4097 4111 4131
rect 4813 4097 4847 4131
rect 4905 4097 4939 4131
rect 5641 4097 5675 4131
rect 6101 4097 6135 4131
rect 6285 4097 6319 4131
rect 6837 4097 6871 4131
rect 7021 4097 7055 4131
rect 7665 4097 7699 4131
rect 9045 4097 9079 4131
rect 5457 3893 5491 3927
rect 6193 3893 6227 3927
rect 9229 3893 9263 3927
rect 3617 3689 3651 3723
rect 4997 3689 5031 3723
rect 6009 3689 6043 3723
rect 9229 3689 9263 3723
rect 4353 3621 4387 3655
rect 3525 3485 3559 3519
rect 3709 3485 3743 3519
rect 4169 3485 4203 3519
rect 4905 3485 4939 3519
rect 6101 3485 6135 3519
rect 7021 3485 7055 3519
rect 7205 3485 7239 3519
rect 8217 3485 8251 3519
rect 9045 3485 9079 3519
rect 7205 3349 7239 3383
rect 8309 3349 8343 3383
rect 4905 3145 4939 3179
rect 6193 3145 6227 3179
rect 7205 3145 7239 3179
rect 7849 3145 7883 3179
rect 9229 3145 9263 3179
rect 4077 3077 4111 3111
rect 3617 3009 3651 3043
rect 4721 3009 4755 3043
rect 4905 3009 4939 3043
rect 5365 3009 5399 3043
rect 5549 3009 5583 3043
rect 6009 3009 6043 3043
rect 7021 3009 7055 3043
rect 7665 3009 7699 3043
rect 8493 3009 8527 3043
rect 8677 3009 8711 3043
rect 9137 3009 9171 3043
rect 9321 3009 9355 3043
rect 5457 2805 5491 2839
rect 8585 2805 8619 2839
rect 3617 2601 3651 2635
rect 4721 2601 4755 2635
rect 8585 2601 8619 2635
rect 6009 2533 6043 2567
rect 9137 2533 9171 2567
rect 3525 2397 3559 2431
rect 3709 2397 3743 2431
rect 4905 2397 4939 2431
rect 5917 2397 5951 2431
rect 6101 2397 6135 2431
rect 6561 2397 6595 2431
rect 6745 2397 6779 2431
rect 7205 2397 7239 2431
rect 7389 2397 7423 2431
rect 8677 2397 8711 2431
rect 9321 2397 9355 2431
rect 6653 2261 6687 2295
rect 7297 2261 7331 2295
rect 3709 2057 3743 2091
rect 4353 2057 4387 2091
rect 5641 2057 5675 2091
rect 6285 2057 6319 2091
rect 7481 2057 7515 2091
rect 9229 2057 9263 2091
rect 3525 1921 3559 1955
rect 4169 1921 4203 1955
rect 4813 1921 4847 1955
rect 4997 1921 5031 1955
rect 5457 1921 5491 1955
rect 6101 1921 6135 1955
rect 6285 1921 6319 1955
rect 6745 1921 6779 1955
rect 6929 1921 6963 1955
rect 7389 1921 7423 1955
rect 9321 1921 9355 1955
rect 8493 1853 8527 1887
rect 8677 1853 8711 1887
rect 4905 1717 4939 1751
rect 6837 1717 6871 1751
rect 3617 1309 3651 1343
rect 3709 1309 3743 1343
rect 4169 1309 4203 1343
rect 4813 1309 4847 1343
rect 5917 1309 5951 1343
rect 6101 1309 6135 1343
rect 6745 1309 6779 1343
rect 7389 1309 7423 1343
rect 6653 1241 6687 1275
rect 4353 1173 4387 1207
rect 4905 1173 4939 1207
rect 6009 1173 6043 1207
rect 7297 1173 7331 1207
<< metal1 >>
rect 1670 15852 1676 15904
rect 1728 15892 1734 15904
rect 2774 15892 2780 15904
rect 1728 15864 2780 15892
rect 1728 15852 1734 15864
rect 2774 15852 2780 15864
rect 2832 15852 2838 15904
rect 920 15802 9844 15824
rect 920 15750 2566 15802
rect 2618 15750 2630 15802
rect 2682 15750 2694 15802
rect 2746 15750 2758 15802
rect 2810 15750 2822 15802
rect 2874 15750 7566 15802
rect 7618 15750 7630 15802
rect 7682 15750 7694 15802
rect 7746 15750 7758 15802
rect 7810 15750 7822 15802
rect 7874 15750 9844 15802
rect 920 15728 9844 15750
rect 2317 15691 2375 15697
rect 2317 15657 2329 15691
rect 2363 15688 2375 15691
rect 2406 15688 2412 15700
rect 2363 15660 2412 15688
rect 2363 15657 2375 15660
rect 2317 15651 2375 15657
rect 2406 15648 2412 15660
rect 2464 15648 2470 15700
rect 5721 15691 5779 15697
rect 5721 15657 5733 15691
rect 5767 15688 5779 15691
rect 6362 15688 6368 15700
rect 5767 15660 6368 15688
rect 5767 15657 5779 15660
rect 5721 15651 5779 15657
rect 6362 15648 6368 15660
rect 6420 15648 6426 15700
rect 4706 15552 4712 15564
rect 2516 15524 4476 15552
rect 4667 15524 4712 15552
rect 1762 15484 1768 15496
rect 1723 15456 1768 15484
rect 1762 15444 1768 15456
rect 1820 15444 1826 15496
rect 2516 15493 2544 15524
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15453 2559 15487
rect 3234 15484 3240 15496
rect 3195 15456 3240 15484
rect 2501 15447 2559 15453
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 2406 15376 2412 15428
rect 2464 15416 2470 15428
rect 2961 15419 3019 15425
rect 2961 15416 2973 15419
rect 2464 15388 2973 15416
rect 2464 15376 2470 15388
rect 2961 15385 2973 15388
rect 3007 15385 3019 15419
rect 2961 15379 3019 15385
rect 3145 15419 3203 15425
rect 3145 15385 3157 15419
rect 3191 15416 3203 15419
rect 4062 15416 4068 15428
rect 3191 15388 4068 15416
rect 3191 15385 3203 15388
rect 3145 15379 3203 15385
rect 4062 15376 4068 15388
rect 4120 15376 4126 15428
rect 4448 15416 4476 15524
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15453 5043 15487
rect 4985 15447 5043 15453
rect 5537 15487 5595 15493
rect 5537 15453 5549 15487
rect 5583 15484 5595 15487
rect 6822 15484 6828 15496
rect 5583 15456 6828 15484
rect 5583 15453 5595 15456
rect 5537 15447 5595 15453
rect 4706 15416 4712 15428
rect 4448 15388 4712 15416
rect 4706 15376 4712 15388
rect 4764 15376 4770 15428
rect 5000 15416 5028 15447
rect 6822 15444 6828 15456
rect 6880 15444 6886 15496
rect 8386 15444 8392 15496
rect 8444 15484 8450 15496
rect 8941 15487 8999 15493
rect 8444 15456 8489 15484
rect 8444 15444 8450 15456
rect 8941 15453 8953 15487
rect 8987 15484 8999 15487
rect 9030 15484 9036 15496
rect 8987 15456 9036 15484
rect 8987 15453 8999 15456
rect 8941 15447 8999 15453
rect 9030 15444 9036 15456
rect 9088 15444 9094 15496
rect 5626 15416 5632 15428
rect 5000 15388 5632 15416
rect 5626 15376 5632 15388
rect 5684 15376 5690 15428
rect 7374 15376 7380 15428
rect 7432 15376 7438 15428
rect 8110 15416 8116 15428
rect 8071 15388 8116 15416
rect 8110 15376 8116 15388
rect 8168 15376 8174 15428
rect 1302 15308 1308 15360
rect 1360 15348 1366 15360
rect 1581 15351 1639 15357
rect 1581 15348 1593 15351
rect 1360 15320 1593 15348
rect 1360 15308 1366 15320
rect 1581 15317 1593 15320
rect 1627 15317 1639 15351
rect 3050 15348 3056 15360
rect 3011 15320 3056 15348
rect 1581 15311 1639 15317
rect 3050 15308 3056 15320
rect 3108 15308 3114 15360
rect 6638 15348 6644 15360
rect 6599 15320 6644 15348
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 9122 15348 9128 15360
rect 9083 15320 9128 15348
rect 9122 15308 9128 15320
rect 9180 15308 9186 15360
rect 920 15258 9844 15280
rect 920 15206 3566 15258
rect 3618 15206 3630 15258
rect 3682 15206 3694 15258
rect 3746 15206 3758 15258
rect 3810 15206 3822 15258
rect 3874 15206 8566 15258
rect 8618 15206 8630 15258
rect 8682 15206 8694 15258
rect 8746 15206 8758 15258
rect 8810 15206 8822 15258
rect 8874 15206 9844 15258
rect 920 15184 9844 15206
rect 5626 15104 5632 15156
rect 5684 15144 5690 15156
rect 6641 15147 6699 15153
rect 6641 15144 6653 15147
rect 5684 15116 6653 15144
rect 5684 15104 5690 15116
rect 6641 15113 6653 15116
rect 6687 15113 6699 15147
rect 6641 15107 6699 15113
rect 1489 15079 1547 15085
rect 1489 15045 1501 15079
rect 1535 15076 1547 15079
rect 1854 15076 1860 15088
rect 1535 15048 1860 15076
rect 1535 15045 1547 15048
rect 1489 15039 1547 15045
rect 1854 15036 1860 15048
rect 1912 15036 1918 15088
rect 2593 15079 2651 15085
rect 2593 15076 2605 15079
rect 2240 15048 2605 15076
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 2240 15008 2268 15048
rect 2593 15045 2605 15048
rect 2639 15076 2651 15079
rect 3421 15079 3479 15085
rect 3421 15076 3433 15079
rect 2639 15048 3433 15076
rect 2639 15045 2651 15048
rect 2593 15039 2651 15045
rect 3421 15045 3433 15048
rect 3467 15076 3479 15079
rect 4154 15076 4160 15088
rect 3467 15048 4160 15076
rect 3467 15045 3479 15048
rect 3421 15039 3479 15045
rect 4154 15036 4160 15048
rect 4212 15036 4218 15088
rect 7374 15036 7380 15088
rect 7432 15036 7438 15088
rect 8113 15079 8171 15085
rect 8113 15045 8125 15079
rect 8159 15076 8171 15079
rect 8202 15076 8208 15088
rect 8159 15048 8208 15076
rect 8159 15045 8171 15048
rect 8113 15039 8171 15045
rect 8202 15036 8208 15048
rect 8260 15036 8266 15088
rect 1719 14980 2268 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 2314 14968 2320 15020
rect 2372 15008 2378 15020
rect 2409 15011 2467 15017
rect 2409 15008 2421 15011
rect 2372 14980 2421 15008
rect 2372 14968 2378 14980
rect 2409 14977 2421 14980
rect 2455 14977 2467 15011
rect 2409 14971 2467 14977
rect 3237 15011 3295 15017
rect 3237 14977 3249 15011
rect 3283 15008 3295 15011
rect 3326 15008 3332 15020
rect 3283 14980 3332 15008
rect 3283 14977 3295 14980
rect 3237 14971 3295 14977
rect 934 14900 940 14952
rect 992 14940 998 14952
rect 2332 14940 2360 14968
rect 3252 14940 3280 14971
rect 3326 14968 3332 14980
rect 3384 14968 3390 15020
rect 4062 15008 4068 15020
rect 4023 14980 4068 15008
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 5718 15008 5724 15020
rect 5679 14980 5724 15008
rect 5718 14968 5724 14980
rect 5776 14968 5782 15020
rect 8938 15008 8944 15020
rect 8899 14980 8944 15008
rect 8938 14968 8944 14980
rect 8996 14968 9002 15020
rect 992 14912 2360 14940
rect 2516 14912 3280 14940
rect 8389 14943 8447 14949
rect 992 14900 998 14912
rect 1394 14832 1400 14884
rect 1452 14872 1458 14884
rect 2516 14872 2544 14912
rect 8389 14909 8401 14943
rect 8435 14940 8447 14943
rect 15930 14940 15936 14952
rect 8435 14912 15936 14940
rect 8435 14909 8447 14912
rect 8389 14903 8447 14909
rect 15930 14900 15936 14912
rect 15988 14900 15994 14952
rect 1452 14844 2544 14872
rect 1452 14832 1458 14844
rect 2774 14832 2780 14884
rect 2832 14872 2838 14884
rect 5169 14875 5227 14881
rect 5169 14872 5181 14875
rect 2832 14844 2877 14872
rect 4172 14844 5181 14872
rect 2832 14832 2838 14844
rect 474 14764 480 14816
rect 532 14804 538 14816
rect 1857 14807 1915 14813
rect 1857 14804 1869 14807
rect 532 14776 1869 14804
rect 532 14764 538 14776
rect 1857 14773 1869 14776
rect 1903 14773 1915 14807
rect 3602 14804 3608 14816
rect 3563 14776 3608 14804
rect 1857 14767 1915 14773
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 4172 14804 4200 14844
rect 5169 14841 5181 14844
rect 5215 14841 5227 14875
rect 5169 14835 5227 14841
rect 4120 14776 4200 14804
rect 4120 14764 4126 14776
rect 4522 14764 4528 14816
rect 4580 14804 4586 14816
rect 4709 14807 4767 14813
rect 4709 14804 4721 14807
rect 4580 14776 4721 14804
rect 4580 14764 4586 14776
rect 4709 14773 4721 14776
rect 4755 14773 4767 14807
rect 4709 14767 4767 14773
rect 9125 14807 9183 14813
rect 9125 14773 9137 14807
rect 9171 14804 9183 14807
rect 11422 14804 11428 14816
rect 9171 14776 11428 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 920 14714 9844 14736
rect 920 14662 2566 14714
rect 2618 14662 2630 14714
rect 2682 14662 2694 14714
rect 2746 14662 2758 14714
rect 2810 14662 2822 14714
rect 2874 14662 7566 14714
rect 7618 14662 7630 14714
rect 7682 14662 7694 14714
rect 7746 14662 7758 14714
rect 7810 14662 7822 14714
rect 7874 14662 9844 14714
rect 13814 14696 13820 14748
rect 13872 14736 13878 14748
rect 16206 14736 16212 14748
rect 13872 14708 16212 14736
rect 13872 14696 13878 14708
rect 16206 14696 16212 14708
rect 16264 14696 16270 14748
rect 920 14640 9844 14662
rect 3970 14492 3976 14544
rect 4028 14492 4034 14544
rect 2961 14467 3019 14473
rect 2961 14433 2973 14467
rect 3007 14464 3019 14467
rect 3988 14464 4016 14492
rect 4798 14464 4804 14476
rect 3007 14436 4016 14464
rect 4759 14436 4804 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 4798 14424 4804 14436
rect 4856 14424 4862 14476
rect 5258 14464 5264 14476
rect 5219 14436 5264 14464
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 6512 14436 8984 14464
rect 6512 14424 6518 14436
rect 3234 14356 3240 14408
rect 3292 14396 3298 14408
rect 3973 14399 4031 14405
rect 3292 14368 3337 14396
rect 3292 14356 3298 14368
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 7745 14399 7803 14405
rect 4019 14368 7512 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 2498 14288 2504 14340
rect 2556 14288 2562 14340
rect 4430 14328 4436 14340
rect 4391 14300 4436 14328
rect 4430 14288 4436 14300
rect 4488 14288 4494 14340
rect 4617 14331 4675 14337
rect 4617 14297 4629 14331
rect 4663 14328 4675 14331
rect 5350 14328 5356 14340
rect 4663 14300 5356 14328
rect 4663 14297 4675 14300
rect 4617 14291 4675 14297
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 3881 14263 3939 14269
rect 3881 14229 3893 14263
rect 3927 14260 3939 14263
rect 3970 14260 3976 14272
rect 3927 14232 3976 14260
rect 3927 14229 3939 14232
rect 3881 14223 3939 14229
rect 3970 14220 3976 14232
rect 4028 14220 4034 14272
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 4632 14260 4660 14291
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 7009 14331 7067 14337
rect 7009 14297 7021 14331
rect 7055 14328 7067 14331
rect 7374 14328 7380 14340
rect 7055 14300 7380 14328
rect 7055 14297 7067 14300
rect 7009 14291 7067 14297
rect 7374 14288 7380 14300
rect 7432 14288 7438 14340
rect 7484 14328 7512 14368
rect 7745 14365 7757 14399
rect 7791 14396 7803 14399
rect 8202 14396 8208 14408
rect 7791 14368 8208 14396
rect 7791 14365 7803 14368
rect 7745 14359 7803 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 8956 14405 8984 14436
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 16022 14464 16028 14476
rect 10744 14436 16028 14464
rect 10744 14424 10750 14436
rect 16022 14424 16028 14436
rect 16080 14424 16086 14476
rect 8941 14399 8999 14405
rect 8941 14365 8953 14399
rect 8987 14396 8999 14399
rect 9490 14396 9496 14408
rect 8987 14368 9496 14396
rect 8987 14365 8999 14368
rect 8941 14359 8999 14365
rect 9490 14356 9496 14368
rect 9548 14356 9554 14408
rect 8386 14328 8392 14340
rect 7484 14300 8392 14328
rect 8386 14288 8392 14300
rect 8444 14288 8450 14340
rect 9125 14331 9183 14337
rect 9125 14297 9137 14331
rect 9171 14328 9183 14331
rect 9398 14328 9404 14340
rect 9171 14300 9404 14328
rect 9171 14297 9183 14300
rect 9125 14291 9183 14297
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 10318 14288 10324 14340
rect 10376 14328 10382 14340
rect 14090 14328 14096 14340
rect 10376 14300 14096 14328
rect 10376 14288 10382 14300
rect 14090 14288 14096 14300
rect 14148 14288 14154 14340
rect 4212 14232 4660 14260
rect 8297 14263 8355 14269
rect 4212 14220 4218 14232
rect 8297 14229 8309 14263
rect 8343 14260 8355 14263
rect 8478 14260 8484 14272
rect 8343 14232 8484 14260
rect 8343 14229 8355 14232
rect 8297 14223 8355 14229
rect 8478 14220 8484 14232
rect 8536 14220 8542 14272
rect 9306 14260 9312 14272
rect 9267 14232 9312 14260
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 920 14170 9844 14192
rect 920 14118 3566 14170
rect 3618 14118 3630 14170
rect 3682 14118 3694 14170
rect 3746 14118 3758 14170
rect 3810 14118 3822 14170
rect 3874 14118 8566 14170
rect 8618 14118 8630 14170
rect 8682 14118 8694 14170
rect 8746 14118 8758 14170
rect 8810 14118 8822 14170
rect 8874 14118 9844 14170
rect 920 14096 9844 14118
rect 2590 14056 2596 14068
rect 2551 14028 2596 14056
rect 2590 14016 2596 14028
rect 2648 14016 2654 14068
rect 5442 14056 5448 14068
rect 5403 14028 5448 14056
rect 5442 14016 5448 14028
rect 5500 14016 5506 14068
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14056 6699 14059
rect 9766 14056 9772 14068
rect 6687 14028 9772 14056
rect 6687 14025 6699 14028
rect 6641 14019 6699 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 2774 13948 2780 14000
rect 2832 13988 2838 14000
rect 2832 13960 3450 13988
rect 2832 13948 2838 13960
rect 7926 13948 7932 14000
rect 7984 13948 7990 14000
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1581 13923 1639 13929
rect 1581 13920 1593 13923
rect 1544 13892 1593 13920
rect 1544 13880 1550 13892
rect 1581 13889 1593 13892
rect 1627 13920 1639 13923
rect 2406 13920 2412 13932
rect 1627 13892 2412 13920
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 3050 13920 3056 13932
rect 3011 13892 3056 13920
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 4522 13920 4528 13932
rect 4483 13892 4528 13920
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 5500 13892 5641 13920
rect 5500 13880 5506 13892
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13889 5871 13923
rect 7098 13920 7104 13932
rect 7059 13892 7104 13920
rect 5813 13883 5871 13889
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 4890 13852 4896 13864
rect 2179 13824 2728 13852
rect 4851 13824 4896 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 2700 13784 2728 13824
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 2958 13784 2964 13796
rect 2700 13756 2964 13784
rect 2958 13744 2964 13756
rect 3016 13744 3022 13796
rect 5074 13744 5080 13796
rect 5132 13784 5138 13796
rect 5828 13784 5856 13883
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 8478 13880 8484 13932
rect 8536 13920 8542 13932
rect 8573 13923 8631 13929
rect 8573 13920 8585 13923
rect 8536 13892 8585 13920
rect 8536 13880 8542 13892
rect 8573 13889 8585 13892
rect 8619 13889 8631 13923
rect 8938 13920 8944 13932
rect 8899 13892 8944 13920
rect 8573 13883 8631 13889
rect 8938 13880 8944 13892
rect 8996 13880 9002 13932
rect 5902 13784 5908 13796
rect 5132 13756 5908 13784
rect 5132 13744 5138 13756
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 2498 13676 2504 13728
rect 2556 13716 2562 13728
rect 3050 13716 3056 13728
rect 2556 13688 3056 13716
rect 2556 13676 2562 13688
rect 3050 13676 3056 13688
rect 3108 13676 3114 13728
rect 920 13626 9844 13648
rect 920 13574 2566 13626
rect 2618 13574 2630 13626
rect 2682 13574 2694 13626
rect 2746 13574 2758 13626
rect 2810 13574 2822 13626
rect 2874 13574 7566 13626
rect 7618 13574 7630 13626
rect 7682 13574 7694 13626
rect 7746 13574 7758 13626
rect 7810 13574 7822 13626
rect 7874 13574 9844 13626
rect 920 13552 9844 13574
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 5442 13376 5448 13388
rect 4479 13348 5448 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 7469 13379 7527 13385
rect 7469 13345 7481 13379
rect 7515 13376 7527 13379
rect 7515 13348 8064 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 3050 13268 3056 13320
rect 3108 13308 3114 13320
rect 3881 13311 3939 13317
rect 3881 13308 3893 13311
rect 3108 13280 3893 13308
rect 3108 13268 3114 13280
rect 3881 13277 3893 13280
rect 3927 13308 3939 13311
rect 3927 13280 5028 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 1486 13240 1492 13252
rect 1447 13212 1492 13240
rect 1486 13200 1492 13212
rect 1544 13200 1550 13252
rect 1578 13132 1584 13184
rect 1636 13172 1642 13184
rect 2777 13175 2835 13181
rect 2777 13172 2789 13175
rect 1636 13144 2789 13172
rect 1636 13132 1642 13144
rect 2777 13141 2789 13144
rect 2823 13141 2835 13175
rect 5000 13172 5028 13280
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 5132 13280 5181 13308
rect 5132 13268 5138 13280
rect 5169 13277 5181 13280
rect 5215 13277 5227 13311
rect 5534 13308 5540 13320
rect 5495 13280 5540 13308
rect 5169 13271 5227 13277
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 8036 13317 8064 13348
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13277 7067 13311
rect 7009 13271 7067 13277
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13277 8079 13311
rect 8021 13271 8079 13277
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13308 8999 13311
rect 9122 13308 9128 13320
rect 8987 13280 9128 13308
rect 8987 13277 8999 13280
rect 8941 13271 8999 13277
rect 6638 13200 6644 13252
rect 6696 13200 6702 13252
rect 7024 13240 7052 13271
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 12158 13240 12164 13252
rect 7024 13212 12164 13240
rect 12158 13200 12164 13212
rect 12216 13200 12222 13252
rect 7282 13172 7288 13184
rect 5000 13144 7288 13172
rect 2777 13135 2835 13141
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 8202 13172 8208 13184
rect 8163 13144 8208 13172
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 9125 13175 9183 13181
rect 9125 13141 9137 13175
rect 9171 13172 9183 13175
rect 15562 13172 15568 13184
rect 9171 13144 15568 13172
rect 9171 13141 9183 13144
rect 9125 13135 9183 13141
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 920 13082 9844 13104
rect 920 13030 3566 13082
rect 3618 13030 3630 13082
rect 3682 13030 3694 13082
rect 3746 13030 3758 13082
rect 3810 13030 3822 13082
rect 3874 13030 8566 13082
rect 8618 13030 8630 13082
rect 8682 13030 8694 13082
rect 8746 13030 8758 13082
rect 8810 13030 8822 13082
rect 8874 13030 9844 13082
rect 13814 13064 13820 13116
rect 13872 13104 13878 13116
rect 15654 13104 15660 13116
rect 13872 13076 15660 13104
rect 13872 13064 13878 13076
rect 15654 13064 15660 13076
rect 15712 13064 15718 13116
rect 920 13008 9844 13030
rect 8294 12968 8300 12980
rect 8255 12940 8300 12968
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 3326 12860 3332 12912
rect 3384 12860 3390 12912
rect 12158 12860 12164 12912
rect 12216 12900 12222 12912
rect 16114 12900 16120 12912
rect 12216 12872 16120 12900
rect 12216 12860 12222 12872
rect 16114 12860 16120 12872
rect 16172 12860 16178 12912
rect 1394 12792 1400 12844
rect 1452 12832 1458 12844
rect 1581 12835 1639 12841
rect 1581 12832 1593 12835
rect 1452 12804 1593 12832
rect 1452 12792 1458 12804
rect 1581 12801 1593 12804
rect 1627 12832 1639 12835
rect 1670 12832 1676 12844
rect 1627 12804 1676 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 2958 12832 2964 12844
rect 2919 12804 2964 12832
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4433 12835 4491 12841
rect 4433 12832 4445 12835
rect 4304 12804 4445 12832
rect 4304 12792 4310 12804
rect 4433 12801 4445 12804
rect 4479 12801 4491 12835
rect 4433 12795 4491 12801
rect 5258 12792 5264 12844
rect 5316 12832 5322 12844
rect 5353 12835 5411 12841
rect 5353 12832 5365 12835
rect 5316 12804 5365 12832
rect 5316 12792 5322 12804
rect 5353 12801 5365 12804
rect 5399 12801 5411 12835
rect 6546 12832 6552 12844
rect 6507 12804 6552 12832
rect 5353 12795 5411 12801
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 9217 12835 9275 12841
rect 7958 12818 9168 12832
rect 7944 12804 9168 12818
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 5629 12767 5687 12773
rect 5629 12733 5641 12767
rect 5675 12764 5687 12767
rect 5810 12764 5816 12776
rect 5675 12736 5816 12764
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 5810 12724 5816 12736
rect 5868 12724 5874 12776
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 6914 12764 6920 12776
rect 6871 12736 6920 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 6914 12724 6920 12736
rect 6972 12724 6978 12776
rect 7282 12724 7288 12776
rect 7340 12764 7346 12776
rect 7944 12764 7972 12804
rect 7340 12736 7972 12764
rect 7340 12724 7346 12736
rect 842 12588 848 12640
rect 900 12628 906 12640
rect 2133 12631 2191 12637
rect 2133 12628 2145 12631
rect 900 12600 2145 12628
rect 900 12588 906 12600
rect 2133 12597 2145 12600
rect 2179 12597 2191 12631
rect 2133 12591 2191 12597
rect 2958 12588 2964 12640
rect 3016 12628 3022 12640
rect 3142 12628 3148 12640
rect 3016 12600 3148 12628
rect 3016 12588 3022 12600
rect 3142 12588 3148 12600
rect 3200 12588 3206 12640
rect 4890 12628 4896 12640
rect 4851 12600 4896 12628
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 9140 12637 9168 12804
rect 9217 12801 9229 12835
rect 9263 12832 9275 12835
rect 15470 12832 15476 12844
rect 9263 12804 15476 12832
rect 9263 12801 9275 12804
rect 9217 12795 9275 12801
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 9125 12631 9183 12637
rect 9125 12597 9137 12631
rect 9171 12628 9183 12631
rect 10134 12628 10140 12640
rect 9171 12600 10140 12628
rect 9171 12597 9183 12600
rect 9125 12591 9183 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 920 12538 9844 12560
rect 920 12486 2566 12538
rect 2618 12486 2630 12538
rect 2682 12486 2694 12538
rect 2746 12486 2758 12538
rect 2810 12486 2822 12538
rect 2874 12486 7566 12538
rect 7618 12486 7630 12538
rect 7682 12486 7694 12538
rect 7746 12486 7758 12538
rect 7810 12486 7822 12538
rect 7874 12486 9844 12538
rect 13170 12520 13176 12572
rect 13228 12560 13234 12572
rect 13906 12560 13912 12572
rect 13228 12532 13912 12560
rect 13228 12520 13234 12532
rect 13906 12520 13912 12532
rect 13964 12520 13970 12572
rect 920 12464 9844 12486
rect 2222 12384 2228 12436
rect 2280 12424 2286 12436
rect 2866 12424 2872 12436
rect 2280 12396 2872 12424
rect 2280 12384 2286 12396
rect 2866 12384 2872 12396
rect 2924 12384 2930 12436
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 15010 12424 15016 12436
rect 6696 12396 15016 12424
rect 6696 12384 6702 12396
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 16482 12424 16488 12436
rect 15344 12396 16488 12424
rect 15344 12384 15350 12396
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 10870 12316 10876 12368
rect 10928 12356 10934 12368
rect 16390 12356 16396 12368
rect 10928 12328 16396 12356
rect 10928 12316 10934 12328
rect 16390 12316 16396 12328
rect 16448 12316 16454 12368
rect 2406 12248 2412 12300
rect 2464 12288 2470 12300
rect 2961 12291 3019 12297
rect 2961 12288 2973 12291
rect 2464 12260 2973 12288
rect 2464 12248 2470 12260
rect 2961 12257 2973 12260
rect 3007 12257 3019 12291
rect 2961 12251 3019 12257
rect 6914 12248 6920 12300
rect 6972 12288 6978 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 6972 12260 7481 12288
rect 6972 12248 6978 12260
rect 7469 12257 7481 12260
rect 7515 12288 7527 12291
rect 8110 12288 8116 12300
rect 7515 12260 8116 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 3234 12180 3240 12232
rect 3292 12220 3298 12232
rect 3789 12223 3847 12229
rect 3292 12192 3337 12220
rect 3292 12180 3298 12192
rect 3789 12189 3801 12223
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12220 4031 12223
rect 4062 12220 4068 12232
rect 4019 12192 4068 12220
rect 4019 12189 4031 12192
rect 3973 12183 4031 12189
rect 3050 12152 3056 12164
rect 2530 12124 3056 12152
rect 3050 12112 3056 12124
rect 3108 12112 3114 12164
rect 3804 12152 3832 12183
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 4433 12223 4491 12229
rect 4433 12220 4445 12223
rect 4304 12192 4445 12220
rect 4304 12180 4310 12192
rect 4433 12189 4445 12192
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 4706 12180 4712 12232
rect 4764 12220 4770 12232
rect 4801 12223 4859 12229
rect 4801 12220 4813 12223
rect 4764 12192 4813 12220
rect 4764 12180 4770 12192
rect 4801 12189 4813 12192
rect 4847 12189 4859 12223
rect 6270 12220 6276 12232
rect 6231 12192 6276 12220
rect 4801 12183 4859 12189
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 8938 12220 8944 12232
rect 8899 12192 8944 12220
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 4338 12152 4344 12164
rect 3804 12124 4344 12152
rect 4338 12112 4344 12124
rect 4396 12112 4402 12164
rect 5902 12112 5908 12164
rect 5960 12112 5966 12164
rect 8478 12112 8484 12164
rect 8536 12152 8542 12164
rect 9125 12155 9183 12161
rect 9125 12152 9137 12155
rect 8536 12124 9137 12152
rect 8536 12112 8542 12124
rect 9125 12121 9137 12124
rect 9171 12152 9183 12155
rect 9398 12152 9404 12164
rect 9171 12124 9404 12152
rect 9171 12121 9183 12124
rect 9125 12115 9183 12121
rect 9398 12112 9404 12124
rect 9456 12112 9462 12164
rect 1489 12087 1547 12093
rect 1489 12053 1501 12087
rect 1535 12084 1547 12087
rect 1670 12084 1676 12096
rect 1535 12056 1676 12084
rect 1535 12053 1547 12056
rect 1489 12047 1547 12053
rect 1670 12044 1676 12056
rect 1728 12044 1734 12096
rect 3881 12087 3939 12093
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 4062 12084 4068 12096
rect 3927 12056 4068 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 6733 12087 6791 12093
rect 6733 12084 6745 12087
rect 5592 12056 6745 12084
rect 5592 12044 5598 12056
rect 6733 12053 6745 12056
rect 6779 12053 6791 12087
rect 6733 12047 6791 12053
rect 8113 12087 8171 12093
rect 8113 12053 8125 12087
rect 8159 12084 8171 12087
rect 8294 12084 8300 12096
rect 8159 12056 8300 12084
rect 8159 12053 8171 12056
rect 8113 12047 8171 12053
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 9309 12087 9367 12093
rect 9309 12053 9321 12087
rect 9355 12084 9367 12087
rect 9950 12084 9956 12096
rect 9355 12056 9956 12084
rect 9355 12053 9367 12056
rect 9309 12047 9367 12053
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 920 11994 9844 12016
rect 920 11942 3566 11994
rect 3618 11942 3630 11994
rect 3682 11942 3694 11994
rect 3746 11942 3758 11994
rect 3810 11942 3822 11994
rect 3874 11942 8566 11994
rect 8618 11942 8630 11994
rect 8682 11942 8694 11994
rect 8746 11942 8758 11994
rect 8810 11942 8822 11994
rect 8874 11942 9844 11994
rect 920 11920 9844 11942
rect 3050 11840 3056 11892
rect 3108 11840 3114 11892
rect 8110 11880 8116 11892
rect 8071 11852 8116 11880
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 9088 11852 9229 11880
rect 9088 11840 9094 11852
rect 9217 11849 9229 11852
rect 9263 11849 9275 11883
rect 9217 11843 9275 11849
rect 11606 11840 11612 11892
rect 11664 11880 11670 11892
rect 16574 11880 16580 11892
rect 11664 11852 16580 11880
rect 11664 11840 11670 11852
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 3068 11812 3096 11840
rect 2898 11784 3096 11812
rect 3234 11772 3240 11824
rect 3292 11812 3298 11824
rect 5810 11812 5816 11824
rect 3292 11784 3648 11812
rect 5771 11784 5816 11812
rect 3292 11772 3298 11784
rect 3620 11753 3648 11784
rect 5810 11772 5816 11784
rect 5868 11772 5874 11824
rect 6546 11812 6552 11824
rect 6380 11784 6552 11812
rect 6380 11753 6408 11784
rect 6546 11772 6552 11784
rect 6604 11772 6610 11824
rect 7282 11772 7288 11824
rect 7340 11772 7346 11824
rect 8846 11812 8852 11824
rect 8807 11784 8852 11812
rect 8846 11772 8852 11784
rect 8904 11772 8910 11824
rect 11422 11772 11428 11824
rect 11480 11812 11486 11824
rect 13722 11812 13728 11824
rect 11480 11784 13728 11812
rect 11480 11772 11486 11784
rect 13722 11772 13728 11784
rect 13780 11772 13786 11824
rect 3605 11747 3663 11753
rect 3605 11713 3617 11747
rect 3651 11744 3663 11747
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 3651 11716 6377 11744
rect 3651 11713 3663 11716
rect 3605 11707 3663 11713
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 8754 11744 8760 11756
rect 8715 11716 8760 11744
rect 6365 11707 6423 11713
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 8938 11704 8944 11756
rect 8996 11744 9002 11756
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8996 11716 9045 11744
rect 8996 11704 9002 11716
rect 9033 11713 9045 11716
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 3234 11636 3240 11688
rect 3292 11676 3298 11688
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 3292 11648 3341 11676
rect 3292 11636 3298 11648
rect 3329 11645 3341 11648
rect 3375 11645 3387 11679
rect 4154 11676 4160 11688
rect 4115 11648 4160 11676
rect 3329 11639 3387 11645
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 6638 11676 6644 11688
rect 6599 11648 6644 11676
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 15470 11568 15476 11620
rect 15528 11608 15534 11620
rect 15746 11608 15752 11620
rect 15528 11580 15752 11608
rect 15528 11568 15534 11580
rect 15746 11568 15752 11580
rect 15804 11568 15810 11620
rect 1854 11540 1860 11552
rect 1815 11512 1860 11540
rect 1854 11500 1860 11512
rect 1912 11500 1918 11552
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 7282 11540 7288 11552
rect 5960 11512 7288 11540
rect 5960 11500 5966 11512
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 7566 11450
rect 7618 11398 7630 11450
rect 7682 11398 7694 11450
rect 7746 11398 7758 11450
rect 7810 11398 7822 11450
rect 7874 11398 9844 11450
rect 920 11376 9844 11398
rect 15286 11364 15292 11416
rect 15344 11404 15350 11416
rect 16666 11404 16672 11416
rect 15344 11376 16672 11404
rect 15344 11364 15350 11376
rect 16666 11364 16672 11376
rect 16724 11364 16730 11416
rect 3237 11339 3295 11345
rect 3237 11305 3249 11339
rect 3283 11336 3295 11339
rect 3326 11336 3332 11348
rect 3283 11308 3332 11336
rect 3283 11305 3295 11308
rect 3237 11299 3295 11305
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 15654 11268 15660 11280
rect 15166 11240 15660 11268
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11200 1639 11203
rect 1762 11200 1768 11212
rect 1627 11172 1768 11200
rect 1627 11169 1639 11172
rect 1581 11163 1639 11169
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 1854 11160 1860 11212
rect 1912 11200 1918 11212
rect 2593 11203 2651 11209
rect 2593 11200 2605 11203
rect 1912 11172 2605 11200
rect 1912 11160 1918 11172
rect 2593 11169 2605 11172
rect 2639 11200 2651 11203
rect 4890 11200 4896 11212
rect 2639 11172 2774 11200
rect 4851 11172 4896 11200
rect 2639 11169 2651 11172
rect 2593 11163 2651 11169
rect 1854 11024 1860 11076
rect 1912 11064 1918 11076
rect 2133 11067 2191 11073
rect 2133 11064 2145 11067
rect 1912 11036 2145 11064
rect 1912 11024 1918 11036
rect 2133 11033 2145 11036
rect 2179 11033 2191 11067
rect 2133 11027 2191 11033
rect 2746 10996 2774 11172
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 5166 11160 5172 11212
rect 5224 11200 5230 11212
rect 8021 11203 8079 11209
rect 8021 11200 8033 11203
rect 5224 11172 8033 11200
rect 5224 11160 5230 11172
rect 8021 11169 8033 11172
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 13354 11160 13360 11212
rect 13412 11200 13418 11212
rect 15166 11200 15194 11240
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 13412 11172 15194 11200
rect 13412 11160 13418 11172
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 7653 11135 7711 11141
rect 7653 11132 7665 11135
rect 7156 11104 7665 11132
rect 7156 11092 7162 11104
rect 7653 11101 7665 11104
rect 7699 11101 7711 11135
rect 7653 11095 7711 11101
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11132 8999 11135
rect 9030 11132 9036 11144
rect 8987 11104 9036 11132
rect 8987 11101 8999 11104
rect 8941 11095 8999 11101
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 11698 11092 11704 11144
rect 11756 11132 11762 11144
rect 13814 11132 13820 11144
rect 11756 11104 13820 11132
rect 11756 11092 11762 11104
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 15470 11092 15476 11144
rect 15528 11132 15534 11144
rect 15654 11132 15660 11144
rect 15528 11104 15660 11132
rect 15528 11092 15534 11104
rect 15654 11092 15660 11104
rect 15712 11092 15718 11144
rect 4154 11024 4160 11076
rect 4212 11064 4218 11076
rect 4249 11067 4307 11073
rect 4249 11064 4261 11067
rect 4212 11036 4261 11064
rect 4212 11024 4218 11036
rect 4249 11033 4261 11036
rect 4295 11033 4307 11067
rect 4249 11027 4307 11033
rect 5442 11024 5448 11076
rect 5500 11064 5506 11076
rect 5537 11067 5595 11073
rect 5537 11064 5549 11067
rect 5500 11036 5549 11064
rect 5500 11024 5506 11036
rect 5537 11033 5549 11036
rect 5583 11033 5595 11067
rect 7190 11064 7196 11076
rect 7151 11036 7196 11064
rect 5537 11027 5595 11033
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 7837 11067 7895 11073
rect 7837 11064 7849 11067
rect 7300 11036 7849 11064
rect 4062 10996 4068 11008
rect 2746 10968 4068 10996
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 5626 10956 5632 11008
rect 5684 10996 5690 11008
rect 7300 10996 7328 11036
rect 7837 11033 7849 11036
rect 7883 11064 7895 11067
rect 8478 11064 8484 11076
rect 7883 11036 8484 11064
rect 7883 11033 7895 11036
rect 7837 11027 7895 11033
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 5684 10968 7328 10996
rect 9125 10999 9183 11005
rect 5684 10956 5690 10968
rect 9125 10965 9137 10999
rect 9171 10996 9183 10999
rect 15470 10996 15476 11008
rect 9171 10968 15476 10996
rect 9171 10965 9183 10968
rect 9125 10959 9183 10965
rect 15470 10956 15476 10968
rect 15528 10956 15534 11008
rect 920 10906 9844 10928
rect 920 10854 3566 10906
rect 3618 10854 3630 10906
rect 3682 10854 3694 10906
rect 3746 10854 3758 10906
rect 3810 10854 3822 10906
rect 3874 10854 8566 10906
rect 8618 10854 8630 10906
rect 8682 10854 8694 10906
rect 8746 10854 8758 10906
rect 8810 10854 8822 10906
rect 8874 10854 9844 10906
rect 15378 10888 15384 10940
rect 15436 10928 15442 10940
rect 15930 10928 15936 10940
rect 15436 10900 15936 10928
rect 15436 10888 15442 10900
rect 15930 10888 15936 10900
rect 15988 10888 15994 10940
rect 920 10832 9844 10854
rect 2314 10752 2320 10804
rect 2372 10792 2378 10804
rect 4801 10795 4859 10801
rect 2372 10764 3188 10792
rect 2372 10752 2378 10764
rect 1394 10724 1400 10736
rect 1355 10696 1400 10724
rect 1394 10684 1400 10696
rect 1452 10684 1458 10736
rect 3160 10724 3188 10764
rect 4801 10761 4813 10795
rect 4847 10792 4859 10795
rect 4890 10792 4896 10804
rect 4847 10764 4896 10792
rect 4847 10761 4859 10764
rect 4801 10755 4859 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 8018 10752 8024 10804
rect 8076 10792 8082 10804
rect 8662 10792 8668 10804
rect 8076 10764 8668 10792
rect 8076 10752 8082 10764
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 9122 10752 9128 10804
rect 9180 10792 9186 10804
rect 15930 10792 15936 10804
rect 9180 10764 15936 10792
rect 9180 10752 9186 10764
rect 15930 10752 15936 10764
rect 15988 10752 15994 10804
rect 5445 10727 5503 10733
rect 3160 10696 3266 10724
rect 5445 10693 5457 10727
rect 5491 10724 5503 10727
rect 5718 10724 5724 10736
rect 5491 10696 5724 10724
rect 5491 10693 5503 10696
rect 5445 10687 5503 10693
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 7190 10684 7196 10736
rect 7248 10684 7254 10736
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10656 1639 10659
rect 2038 10656 2044 10668
rect 1627 10628 2044 10656
rect 1627 10625 1639 10628
rect 1581 10619 1639 10625
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2130 10616 2136 10668
rect 2188 10656 2194 10668
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2188 10628 2881 10656
rect 2188 10616 2194 10628
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4614 10656 4620 10668
rect 4387 10628 4620 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 5626 10656 5632 10668
rect 5408 10628 5632 10656
rect 5408 10616 5414 10628
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 6178 10616 6184 10668
rect 6236 10656 6242 10668
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6236 10628 6837 10656
rect 6236 10616 6242 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 8294 10656 8300 10668
rect 8255 10628 8300 10656
rect 6825 10619 6883 10625
rect 8294 10616 8300 10628
rect 8352 10616 8358 10668
rect 8386 10616 8392 10668
rect 8444 10656 8450 10668
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 8444 10628 9137 10656
rect 8444 10616 8450 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 2498 10588 2504 10600
rect 2459 10560 2504 10588
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 7926 10548 7932 10600
rect 7984 10588 7990 10600
rect 8665 10591 8723 10597
rect 7984 10560 8616 10588
rect 7984 10548 7990 10560
rect 8588 10520 8616 10560
rect 8665 10557 8677 10591
rect 8711 10588 8723 10591
rect 9217 10591 9275 10597
rect 9217 10588 9229 10591
rect 8711 10560 9229 10588
rect 8711 10557 8723 10560
rect 8665 10551 8723 10557
rect 9217 10557 9229 10560
rect 9263 10557 9275 10591
rect 9217 10551 9275 10557
rect 16298 10520 16304 10532
rect 8588 10492 16304 10520
rect 16298 10480 16304 10492
rect 16356 10480 16362 10532
rect 1765 10455 1823 10461
rect 1765 10421 1777 10455
rect 1811 10452 1823 10455
rect 5258 10452 5264 10464
rect 1811 10424 5264 10452
rect 1811 10421 1823 10424
rect 1765 10415 1823 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5810 10452 5816 10464
rect 5771 10424 5816 10452
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 6086 10412 6092 10464
rect 6144 10452 6150 10464
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 6144 10424 6377 10452
rect 6144 10412 6150 10424
rect 6365 10421 6377 10424
rect 6411 10421 6423 10455
rect 6365 10415 6423 10421
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 7566 10362
rect 7618 10310 7630 10362
rect 7682 10310 7694 10362
rect 7746 10310 7758 10362
rect 7810 10310 7822 10362
rect 7874 10310 9844 10362
rect 920 10288 9844 10310
rect 2130 10248 2136 10260
rect 2091 10220 2136 10248
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 8938 10248 8944 10260
rect 8899 10220 8944 10248
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9122 10248 9128 10260
rect 9083 10220 9128 10248
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 16758 10248 16764 10260
rect 10192 10220 16764 10248
rect 10192 10208 10198 10220
rect 16758 10208 16764 10220
rect 16816 10208 16822 10260
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 1670 10112 1676 10124
rect 1627 10084 1676 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 2222 10072 2228 10124
rect 2280 10112 2286 10124
rect 2593 10115 2651 10121
rect 2593 10112 2605 10115
rect 2280 10084 2605 10112
rect 2280 10072 2286 10084
rect 2593 10081 2605 10084
rect 2639 10081 2651 10115
rect 4062 10112 4068 10124
rect 4023 10084 4068 10112
rect 2593 10075 2651 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10112 8355 10115
rect 9398 10112 9404 10124
rect 8343 10084 9404 10112
rect 8343 10081 8355 10084
rect 8297 10075 8355 10081
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 3418 10004 3424 10056
rect 3476 10044 3482 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3476 10016 3801 10044
rect 3476 10004 3482 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 5994 10044 6000 10056
rect 5955 10016 6000 10044
rect 3789 10007 3847 10013
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6362 10044 6368 10056
rect 6323 10016 6368 10044
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 8478 10044 8484 10056
rect 7883 10016 8484 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 5902 9976 5908 9988
rect 5290 9948 5908 9976
rect 5902 9936 5908 9948
rect 5960 9936 5966 9988
rect 6914 9936 6920 9988
rect 6972 9936 6978 9988
rect 8202 9936 8208 9988
rect 8260 9976 8266 9988
rect 9309 9979 9367 9985
rect 9309 9976 9321 9979
rect 8260 9948 9321 9976
rect 8260 9936 8266 9948
rect 9309 9945 9321 9948
rect 9355 9945 9367 9979
rect 9309 9939 9367 9945
rect 3234 9908 3240 9920
rect 3195 9880 3240 9908
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 5537 9911 5595 9917
rect 5537 9877 5549 9911
rect 5583 9908 5595 9911
rect 6638 9908 6644 9920
rect 5583 9880 6644 9908
rect 5583 9877 5595 9880
rect 5537 9871 5595 9877
rect 6638 9868 6644 9880
rect 6696 9908 6702 9920
rect 6822 9908 6828 9920
rect 6696 9880 6828 9908
rect 6696 9868 6702 9880
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 8018 9908 8024 9920
rect 7979 9880 8024 9908
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 9122 9917 9128 9920
rect 9109 9911 9128 9917
rect 9109 9908 9121 9911
rect 8720 9880 9121 9908
rect 8720 9868 8726 9880
rect 9109 9877 9121 9880
rect 9109 9871 9128 9877
rect 9122 9868 9128 9871
rect 9180 9868 9186 9920
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 15102 9908 15108 9920
rect 13872 9880 15108 9908
rect 13872 9868 13878 9880
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 16206 9840 16212 9852
rect 920 9818 9844 9840
rect 920 9766 3566 9818
rect 3618 9766 3630 9818
rect 3682 9766 3694 9818
rect 3746 9766 3758 9818
rect 3810 9766 3822 9818
rect 3874 9766 8566 9818
rect 8618 9766 8630 9818
rect 8682 9766 8694 9818
rect 8746 9766 8758 9818
rect 8810 9766 8822 9818
rect 8874 9766 9844 9818
rect 920 9744 9844 9766
rect 11624 9812 16212 9840
rect 11624 9704 11652 9812
rect 16206 9800 16212 9812
rect 16264 9800 16270 9852
rect 11698 9732 11704 9784
rect 11756 9772 11762 9784
rect 16850 9772 16856 9784
rect 11756 9744 16856 9772
rect 11756 9732 11762 9744
rect 16850 9732 16856 9744
rect 16908 9732 16914 9784
rect 9140 9676 11652 9704
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 3234 9636 3240 9648
rect 3016 9608 3240 9636
rect 3016 9596 3022 9608
rect 3234 9596 3240 9608
rect 3292 9596 3298 9648
rect 4338 9596 4344 9648
rect 4396 9596 4402 9648
rect 7374 9636 7380 9648
rect 7335 9608 7380 9636
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 9140 9645 9168 9676
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 15102 9704 15108 9716
rect 13872 9676 15108 9704
rect 13872 9664 13878 9676
rect 15102 9664 15108 9676
rect 15160 9664 15166 9716
rect 9125 9639 9183 9645
rect 9125 9605 9137 9639
rect 9171 9605 9183 9639
rect 9125 9599 9183 9605
rect 3050 9568 3056 9580
rect 3011 9540 3056 9568
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9568 3571 9571
rect 3970 9568 3976 9580
rect 3559 9540 3976 9568
rect 3559 9537 3571 9540
rect 3513 9531 3571 9537
rect 3970 9528 3976 9540
rect 4028 9528 4034 9580
rect 5350 9568 5356 9580
rect 5311 9540 5356 9568
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 6457 9571 6515 9577
rect 6457 9537 6469 9571
rect 6503 9568 6515 9571
rect 7006 9568 7012 9580
rect 6503 9540 7012 9568
rect 6503 9537 6515 9540
rect 6457 9531 6515 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 15194 9528 15200 9580
rect 15252 9568 15258 9580
rect 15470 9568 15476 9580
rect 15252 9540 15476 9568
rect 15252 9528 15258 9540
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 16850 9568 16856 9580
rect 16540 9540 16856 9568
rect 16540 9528 16546 9540
rect 16850 9528 16856 9540
rect 16908 9528 16914 9580
rect 1489 9503 1547 9509
rect 1489 9469 1501 9503
rect 1535 9500 1547 9503
rect 2222 9500 2228 9512
rect 1535 9472 2228 9500
rect 1535 9469 1547 9472
rect 1489 9463 1547 9469
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 2682 9500 2688 9512
rect 2643 9472 2688 9500
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3016 9472 3893 9500
rect 3016 9460 3022 9472
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 5810 9500 5816 9512
rect 5771 9472 5816 9500
rect 3881 9463 3939 9469
rect 5810 9460 5816 9472
rect 5868 9460 5874 9512
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 4856 9336 6561 9364
rect 4856 9324 4862 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 6917 9367 6975 9373
rect 6917 9333 6929 9367
rect 6963 9364 6975 9367
rect 9030 9364 9036 9376
rect 6963 9336 9036 9364
rect 6963 9333 6975 9336
rect 6917 9327 6975 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 7566 9274
rect 7618 9222 7630 9274
rect 7682 9222 7694 9274
rect 7746 9222 7758 9274
rect 7810 9222 7822 9274
rect 7874 9222 9844 9274
rect 920 9200 9844 9222
rect 13814 9188 13820 9240
rect 13872 9228 13878 9240
rect 15562 9228 15568 9240
rect 13872 9200 15568 9228
rect 13872 9188 13878 9200
rect 15562 9188 15568 9200
rect 15620 9188 15626 9240
rect 4706 9160 4712 9172
rect 4667 9132 4712 9160
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 1762 9024 1768 9036
rect 1723 8996 1768 9024
rect 1762 8984 1768 8996
rect 1820 8984 1826 9036
rect 3050 8984 3056 9036
rect 3108 9024 3114 9036
rect 3326 9024 3332 9036
rect 3108 8996 3332 9024
rect 3108 8984 3114 8996
rect 3326 8984 3332 8996
rect 3384 9024 3390 9036
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 3384 8996 4077 9024
rect 3384 8984 3390 8996
rect 4065 8993 4077 8996
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 7653 9027 7711 9033
rect 7653 9024 7665 9027
rect 7064 8996 7665 9024
rect 7064 8984 7070 8996
rect 7653 8993 7665 8996
rect 7699 8993 7711 9027
rect 7653 8987 7711 8993
rect 1486 8956 1492 8968
rect 1447 8928 1492 8956
rect 1486 8916 1492 8928
rect 1544 8916 1550 8968
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 5261 8959 5319 8965
rect 5261 8956 5273 8959
rect 4212 8928 5273 8956
rect 4212 8916 4218 8928
rect 5261 8925 5273 8928
rect 5307 8956 5319 8959
rect 5442 8956 5448 8968
rect 5307 8928 5448 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 7282 8916 7288 8968
rect 7340 8956 7346 8968
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 7340 8928 7481 8956
rect 7340 8916 7346 8928
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 9030 8956 9036 8968
rect 8991 8928 9036 8956
rect 7469 8919 7527 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 3326 8888 3332 8900
rect 2990 8860 3332 8888
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 1762 8780 1768 8832
rect 1820 8820 1826 8832
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 1820 8792 3249 8820
rect 1820 8780 1826 8792
rect 3237 8789 3249 8792
rect 3283 8789 3295 8823
rect 6546 8820 6552 8832
rect 6507 8792 6552 8820
rect 3237 8783 3295 8789
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 9122 8820 9128 8832
rect 9083 8792 9128 8820
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 15286 8820 15292 8832
rect 9640 8792 15292 8820
rect 9640 8780 9646 8792
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 920 8730 9844 8752
rect 920 8678 3566 8730
rect 3618 8678 3630 8730
rect 3682 8678 3694 8730
rect 3746 8678 3758 8730
rect 3810 8678 3822 8730
rect 3874 8678 8566 8730
rect 8618 8678 8630 8730
rect 8682 8678 8694 8730
rect 8746 8678 8758 8730
rect 8810 8678 8822 8730
rect 8874 8678 9844 8730
rect 920 8656 9844 8678
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 4856 8588 5089 8616
rect 4856 8576 4862 8588
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 5626 8616 5632 8628
rect 5587 8588 5632 8616
rect 5077 8579 5135 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 6362 8616 6368 8628
rect 6323 8588 6368 8616
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 16482 8616 16488 8628
rect 9548 8588 16488 8616
rect 9548 8576 9554 8588
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 3878 8508 3884 8560
rect 3936 8508 3942 8560
rect 9122 8548 9128 8560
rect 9083 8520 9128 8548
rect 9122 8508 9128 8520
rect 9180 8508 9186 8560
rect 1762 8480 1768 8492
rect 1723 8452 1768 8480
rect 1762 8440 1768 8452
rect 1820 8440 1826 8492
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 3145 8483 3203 8489
rect 3145 8480 3157 8483
rect 2363 8452 3157 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 3145 8449 3157 8452
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 4430 8440 4436 8492
rect 4488 8480 4494 8492
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 4488 8452 4629 8480
rect 4488 8440 4494 8452
rect 4617 8449 4629 8452
rect 4663 8449 4675 8483
rect 5810 8480 5816 8492
rect 5771 8452 5816 8480
rect 4617 8443 4675 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 6914 8480 6920 8492
rect 6875 8452 6920 8480
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8480 9367 8483
rect 9582 8480 9588 8492
rect 9355 8452 9588 8480
rect 9355 8449 9367 8452
rect 9309 8443 9367 8449
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 8202 8412 8208 8424
rect 2832 8384 2877 8412
rect 8163 8384 8208 8412
rect 2832 8372 2838 8384
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 10502 8372 10508 8424
rect 10560 8412 10566 8424
rect 15746 8412 15752 8424
rect 10560 8384 15752 8412
rect 10560 8372 10566 8384
rect 15746 8372 15752 8384
rect 15804 8372 15810 8424
rect 6454 8304 6460 8356
rect 6512 8344 6518 8356
rect 7006 8344 7012 8356
rect 6512 8316 7012 8344
rect 6512 8304 6518 8316
rect 7006 8304 7012 8316
rect 7064 8304 7070 8356
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 7566 8186
rect 7618 8134 7630 8186
rect 7682 8134 7694 8186
rect 7746 8134 7758 8186
rect 7810 8134 7822 8186
rect 7874 8134 9844 8186
rect 920 8112 9844 8134
rect 5258 8032 5264 8084
rect 5316 8072 5322 8084
rect 9490 8072 9496 8084
rect 5316 8044 9496 8072
rect 5316 8032 5322 8044
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 3234 7896 3240 7948
rect 3292 7936 3298 7948
rect 3789 7939 3847 7945
rect 3789 7936 3801 7939
rect 3292 7908 3801 7936
rect 3292 7896 3298 7908
rect 3789 7905 3801 7908
rect 3835 7905 3847 7939
rect 3789 7899 3847 7905
rect 1489 7871 1547 7877
rect 1489 7837 1501 7871
rect 1535 7868 1547 7871
rect 1578 7868 1584 7880
rect 1535 7840 1584 7868
rect 1535 7837 1547 7840
rect 1489 7831 1547 7837
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7374 7868 7380 7880
rect 7055 7840 7380 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 8018 7868 8024 7880
rect 7979 7840 8024 7868
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 9088 7840 9137 7868
rect 9088 7828 9094 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 3234 7800 3240 7812
rect 3195 7772 3240 7800
rect 3234 7760 3240 7772
rect 3292 7760 3298 7812
rect 5258 7800 5264 7812
rect 5219 7772 5264 7800
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 8941 7803 8999 7809
rect 8941 7800 8953 7803
rect 8168 7772 8953 7800
rect 8168 7760 8174 7772
rect 8941 7769 8953 7772
rect 8987 7800 8999 7803
rect 8987 7772 9168 7800
rect 8987 7769 8999 7772
rect 8941 7763 8999 7769
rect 9140 7744 9168 7772
rect 4433 7735 4491 7741
rect 4433 7701 4445 7735
rect 4479 7732 4491 7735
rect 4982 7732 4988 7744
rect 4479 7704 4988 7732
rect 4479 7701 4491 7704
rect 4433 7695 4491 7701
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7469 7735 7527 7741
rect 7469 7732 7481 7735
rect 7064 7704 7481 7732
rect 7064 7692 7070 7704
rect 7469 7701 7481 7704
rect 7515 7701 7527 7735
rect 7469 7695 7527 7701
rect 9122 7692 9128 7744
rect 9180 7692 9186 7744
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 9309 7735 9367 7741
rect 9309 7732 9321 7735
rect 9272 7704 9321 7732
rect 9272 7692 9278 7704
rect 9309 7701 9321 7704
rect 9355 7701 9367 7735
rect 9309 7695 9367 7701
rect 920 7642 9844 7664
rect 920 7590 3566 7642
rect 3618 7590 3630 7642
rect 3682 7590 3694 7642
rect 3746 7590 3758 7642
rect 3810 7590 3822 7642
rect 3874 7590 8566 7642
rect 8618 7590 8630 7642
rect 8682 7590 8694 7642
rect 8746 7590 8758 7642
rect 8810 7590 8822 7642
rect 8874 7590 9844 7642
rect 920 7568 9844 7590
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 5408 7500 5825 7528
rect 5408 7488 5414 7500
rect 5813 7497 5825 7500
rect 5859 7528 5871 7531
rect 8018 7528 8024 7540
rect 5859 7500 8024 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 8938 7488 8944 7540
rect 8996 7528 9002 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8996 7500 9137 7528
rect 8996 7488 9002 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9125 7491 9183 7497
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 1857 7463 1915 7469
rect 1857 7460 1869 7463
rect 1544 7432 1869 7460
rect 1544 7420 1550 7432
rect 1857 7429 1869 7432
rect 1903 7460 1915 7463
rect 3418 7460 3424 7472
rect 1903 7432 3424 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 3418 7420 3424 7432
rect 3476 7420 3482 7472
rect 3605 7463 3663 7469
rect 3605 7429 3617 7463
rect 3651 7460 3663 7463
rect 4062 7460 4068 7472
rect 3651 7432 4068 7460
rect 3651 7429 3663 7432
rect 3605 7423 3663 7429
rect 4062 7420 4068 7432
rect 4120 7420 4126 7472
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 4341 7463 4399 7469
rect 4341 7460 4353 7463
rect 4304 7432 4353 7460
rect 4304 7420 4310 7432
rect 4341 7429 4353 7432
rect 4387 7429 4399 7463
rect 4341 7423 4399 7429
rect 4798 7420 4804 7472
rect 4856 7420 4862 7472
rect 7098 7420 7104 7472
rect 7156 7420 7162 7472
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 8076 7364 8217 7392
rect 8076 7352 8082 7364
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 9490 7392 9496 7404
rect 9355 7364 9496 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 3418 7284 3424 7336
rect 3476 7324 3482 7336
rect 4065 7327 4123 7333
rect 4065 7324 4077 7327
rect 3476 7296 4077 7324
rect 3476 7284 3482 7296
rect 4065 7293 4077 7296
rect 4111 7293 4123 7327
rect 6362 7324 6368 7336
rect 6323 7296 6368 7324
rect 4065 7287 4123 7293
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 6733 7327 6791 7333
rect 6733 7293 6745 7327
rect 6779 7324 6791 7327
rect 6914 7324 6920 7336
rect 6779 7296 6920 7324
rect 6779 7293 6791 7296
rect 6733 7287 6791 7293
rect 6914 7284 6920 7296
rect 6972 7284 6978 7336
rect 8665 7191 8723 7197
rect 8665 7157 8677 7191
rect 8711 7188 8723 7191
rect 8938 7188 8944 7200
rect 8711 7160 8944 7188
rect 8711 7157 8723 7160
rect 8665 7151 8723 7157
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 7566 7098
rect 7618 7046 7630 7098
rect 7682 7046 7694 7098
rect 7746 7046 7758 7098
rect 7810 7046 7822 7098
rect 7874 7046 9844 7098
rect 10778 7080 10784 7132
rect 10836 7120 10842 7132
rect 15378 7120 15384 7132
rect 10836 7092 15384 7120
rect 10836 7080 10842 7092
rect 15378 7080 15384 7092
rect 15436 7080 15442 7132
rect 920 7024 9844 7046
rect 10870 6944 10876 6996
rect 10928 6984 10934 6996
rect 16942 6984 16948 6996
rect 10928 6956 16948 6984
rect 10928 6944 10934 6956
rect 16942 6944 16948 6956
rect 17000 6944 17006 6996
rect 4246 6916 4252 6928
rect 4080 6888 4252 6916
rect 1486 6848 1492 6860
rect 1447 6820 1492 6848
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 1762 6848 1768 6860
rect 1723 6820 1768 6848
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 4080 6848 4108 6888
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 3927 6820 4108 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 4798 6848 4804 6860
rect 4212 6820 4804 6848
rect 4212 6808 4218 6820
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 16022 6848 16028 6860
rect 11204 6820 16028 6848
rect 11204 6808 11210 6820
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 3326 6780 3332 6792
rect 2898 6752 3332 6780
rect 3326 6740 3332 6752
rect 3384 6780 3390 6792
rect 4172 6780 4200 6808
rect 3384 6752 4278 6780
rect 3384 6740 3390 6752
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 6086 6780 6092 6792
rect 5684 6752 5729 6780
rect 6047 6752 6092 6780
rect 5684 6740 5690 6752
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 6454 6780 6460 6792
rect 6415 6752 6460 6780
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7524 6752 7941 6780
rect 7524 6740 7530 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8168 6752 8953 6780
rect 8168 6740 8174 6752
rect 8941 6749 8953 6752
rect 8987 6780 8999 6783
rect 9306 6780 9312 6792
rect 8987 6752 9312 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 5353 6715 5411 6721
rect 5353 6681 5365 6715
rect 5399 6712 5411 6715
rect 5399 6684 5580 6712
rect 5399 6681 5411 6684
rect 5353 6675 5411 6681
rect 5552 6656 5580 6684
rect 7098 6672 7104 6724
rect 7156 6672 7162 6724
rect 8846 6712 8852 6724
rect 7944 6684 8852 6712
rect 7944 6656 7972 6684
rect 8846 6672 8852 6684
rect 8904 6712 8910 6724
rect 9125 6715 9183 6721
rect 9125 6712 9137 6715
rect 8904 6684 9137 6712
rect 8904 6672 8910 6684
rect 9125 6681 9137 6684
rect 9171 6681 9183 6715
rect 9125 6675 9183 6681
rect 13170 6672 13176 6724
rect 13228 6712 13234 6724
rect 13630 6712 13636 6724
rect 13228 6684 13636 6712
rect 13228 6672 13234 6684
rect 13630 6672 13636 6684
rect 13688 6672 13694 6724
rect 3237 6647 3295 6653
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 3326 6644 3332 6656
rect 3283 6616 3332 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 5534 6604 5540 6656
rect 5592 6604 5598 6656
rect 7926 6604 7932 6656
rect 7984 6604 7990 6656
rect 8389 6647 8447 6653
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 9030 6644 9036 6656
rect 8435 6616 9036 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 9306 6644 9312 6656
rect 9267 6616 9312 6644
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 920 6554 9844 6576
rect 920 6502 3566 6554
rect 3618 6502 3630 6554
rect 3682 6502 3694 6554
rect 3746 6502 3758 6554
rect 3810 6502 3822 6554
rect 3874 6502 8566 6554
rect 8618 6502 8630 6554
rect 8682 6502 8694 6554
rect 8746 6502 8758 6554
rect 8810 6502 8822 6554
rect 8874 6502 9844 6554
rect 920 6480 9844 6502
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 2958 6440 2964 6452
rect 2363 6412 2964 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 3237 6443 3295 6449
rect 3237 6440 3249 6443
rect 3108 6412 3249 6440
rect 3108 6400 3114 6412
rect 3237 6409 3249 6412
rect 3283 6409 3295 6443
rect 3237 6403 3295 6409
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 5626 6440 5632 6452
rect 3476 6412 5632 6440
rect 3476 6400 3482 6412
rect 4154 6332 4160 6384
rect 4212 6332 4218 6384
rect 5000 6313 5028 6412
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 15654 6440 15660 6452
rect 13872 6412 15660 6440
rect 13872 6400 13878 6412
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 7374 6332 7380 6384
rect 7432 6332 7438 6384
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 5994 6304 6000 6316
rect 5859 6276 6000 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 7006 6304 7012 6316
rect 6963 6276 7012 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6304 8447 6307
rect 9766 6304 9772 6316
rect 8435 6276 9772 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 1765 6239 1823 6245
rect 1765 6205 1777 6239
rect 1811 6236 1823 6239
rect 3326 6236 3332 6248
rect 1811 6208 3332 6236
rect 1811 6205 1823 6208
rect 1765 6199 1823 6205
rect 3326 6196 3332 6208
rect 3384 6196 3390 6248
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 5350 6236 5356 6248
rect 4755 6208 5356 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 6549 6239 6607 6245
rect 6549 6205 6561 6239
rect 6595 6236 6607 6239
rect 6822 6236 6828 6248
rect 6595 6208 6828 6236
rect 6595 6205 6607 6208
rect 6549 6199 6607 6205
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 13078 6196 13084 6248
rect 13136 6236 13142 6248
rect 16850 6236 16856 6248
rect 13136 6208 16856 6236
rect 13136 6196 13142 6208
rect 16850 6196 16856 6208
rect 16908 6196 16914 6248
rect 5629 6171 5687 6177
rect 5629 6137 5641 6171
rect 5675 6168 5687 6171
rect 5718 6168 5724 6180
rect 5675 6140 5724 6168
rect 5675 6137 5687 6140
rect 5629 6131 5687 6137
rect 5718 6128 5724 6140
rect 5776 6128 5782 6180
rect 13814 6128 13820 6180
rect 13872 6168 13878 6180
rect 15930 6168 15936 6180
rect 13872 6140 15936 6168
rect 13872 6128 13878 6140
rect 15930 6128 15936 6140
rect 15988 6128 15994 6180
rect 8846 6100 8852 6112
rect 8807 6072 8852 6100
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 7566 6010
rect 7618 5958 7630 6010
rect 7682 5958 7694 6010
rect 7746 5958 7758 6010
rect 7810 5958 7822 6010
rect 7874 5958 9844 6010
rect 920 5936 9844 5958
rect 2406 5856 2412 5908
rect 2464 5896 2470 5908
rect 2501 5899 2559 5905
rect 2501 5896 2513 5899
rect 2464 5868 2513 5896
rect 2464 5856 2470 5868
rect 2501 5865 2513 5868
rect 2547 5865 2559 5899
rect 5534 5896 5540 5908
rect 5495 5868 5540 5896
rect 2501 5859 2559 5865
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 6972 5868 7021 5896
rect 6972 5856 6978 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 8294 5896 8300 5908
rect 8255 5868 8300 5896
rect 7009 5859 7067 5865
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 1765 5831 1823 5837
rect 1765 5797 1777 5831
rect 1811 5828 1823 5831
rect 2682 5828 2688 5840
rect 1811 5800 2688 5828
rect 1811 5797 1823 5800
rect 1765 5791 1823 5797
rect 2682 5788 2688 5800
rect 2740 5788 2746 5840
rect 3418 5720 3424 5772
rect 3476 5760 3482 5772
rect 3789 5763 3847 5769
rect 3789 5760 3801 5763
rect 3476 5732 3801 5760
rect 3476 5720 3482 5732
rect 3789 5729 3801 5732
rect 3835 5729 3847 5763
rect 5552 5760 5580 5856
rect 6365 5763 6423 5769
rect 6365 5760 6377 5763
rect 5552 5732 6377 5760
rect 3789 5723 3847 5729
rect 6365 5729 6377 5732
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 8294 5720 8300 5772
rect 8352 5760 8358 5772
rect 9122 5760 9128 5772
rect 8352 5732 9128 5760
rect 8352 5720 8358 5732
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 1946 5692 1952 5704
rect 1907 5664 1952 5692
rect 1946 5652 1952 5664
rect 2004 5652 2010 5704
rect 2314 5652 2320 5704
rect 2372 5692 2378 5704
rect 2685 5695 2743 5701
rect 2685 5692 2697 5695
rect 2372 5664 2697 5692
rect 2372 5652 2378 5664
rect 2685 5661 2697 5664
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5692 7803 5695
rect 8202 5692 8208 5704
rect 7791 5664 8208 5692
rect 7791 5661 7803 5664
rect 7745 5655 7803 5661
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 9214 5692 9220 5704
rect 9175 5664 9220 5692
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 3326 5584 3332 5636
rect 3384 5624 3390 5636
rect 4065 5627 4123 5633
rect 4065 5624 4077 5627
rect 3384 5596 4077 5624
rect 3384 5584 3390 5596
rect 4065 5593 4077 5596
rect 4111 5593 4123 5627
rect 4065 5587 4123 5593
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 4212 5596 4554 5624
rect 4212 5584 4218 5596
rect 4448 5556 4476 5596
rect 5994 5584 6000 5636
rect 6052 5624 6058 5636
rect 8941 5627 8999 5633
rect 8941 5624 8953 5627
rect 6052 5596 8953 5624
rect 6052 5584 6058 5596
rect 8404 5568 8432 5596
rect 8941 5593 8953 5596
rect 8987 5593 8999 5627
rect 8941 5587 8999 5593
rect 9125 5627 9183 5633
rect 9125 5593 9137 5627
rect 9171 5624 9183 5627
rect 9490 5624 9496 5636
rect 9171 5596 9496 5624
rect 9171 5593 9183 5596
rect 9125 5587 9183 5593
rect 9490 5584 9496 5596
rect 9548 5624 9554 5636
rect 13814 5624 13820 5636
rect 9548 5596 13820 5624
rect 9548 5584 9554 5596
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 5534 5556 5540 5568
rect 4448 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 7561 5559 7619 5565
rect 7561 5556 7573 5559
rect 6604 5528 7573 5556
rect 6604 5516 6610 5528
rect 7561 5525 7573 5528
rect 7607 5556 7619 5559
rect 7926 5556 7932 5568
rect 7607 5528 7932 5556
rect 7607 5525 7619 5528
rect 7561 5519 7619 5525
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 8386 5516 8392 5568
rect 8444 5516 8450 5568
rect 9030 5556 9036 5568
rect 8991 5528 9036 5556
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 920 5466 9844 5488
rect 920 5414 3566 5466
rect 3618 5414 3630 5466
rect 3682 5414 3694 5466
rect 3746 5414 3758 5466
rect 3810 5414 3822 5466
rect 3874 5414 8566 5466
rect 8618 5414 8630 5466
rect 8682 5414 8694 5466
rect 8746 5414 8758 5466
rect 8810 5414 8822 5466
rect 8874 5414 9844 5466
rect 920 5392 9844 5414
rect 106 5312 112 5364
rect 164 5352 170 5364
rect 2406 5352 2412 5364
rect 164 5324 2412 5352
rect 164 5312 170 5324
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 4062 5352 4068 5364
rect 4023 5324 4068 5352
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 5813 5355 5871 5361
rect 5813 5321 5825 5355
rect 5859 5352 5871 5355
rect 6454 5352 6460 5364
rect 5859 5324 6460 5352
rect 5859 5321 5871 5324
rect 5813 5315 5871 5321
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 7285 5355 7343 5361
rect 7285 5352 7297 5355
rect 6972 5324 7297 5352
rect 6972 5312 6978 5324
rect 7285 5321 7297 5324
rect 7331 5321 7343 5355
rect 7285 5315 7343 5321
rect 6730 5284 6736 5296
rect 5276 5256 6736 5284
rect 5276 5228 5304 5256
rect 6730 5244 6736 5256
rect 6788 5284 6794 5296
rect 9214 5284 9220 5296
rect 6788 5256 7236 5284
rect 9175 5256 9220 5284
rect 6788 5244 6794 5256
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 5258 5216 5264 5228
rect 4203 5188 5264 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 5868 5188 6377 5216
rect 5868 5176 5874 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6546 5176 6552 5228
rect 6604 5216 6610 5228
rect 7208 5225 7236 5256
rect 9214 5244 9220 5256
rect 9272 5244 9278 5296
rect 7193 5219 7251 5225
rect 6604 5188 6697 5216
rect 6604 5176 6610 5188
rect 7193 5185 7205 5219
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 7926 5176 7932 5228
rect 7984 5216 7990 5228
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 7984 5188 9137 5216
rect 7984 5176 7990 5188
rect 9125 5185 9137 5188
rect 9171 5216 9183 5219
rect 10042 5216 10048 5228
rect 9171 5188 10048 5216
rect 9171 5185 9183 5188
rect 9125 5179 9183 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 5169 5151 5227 5157
rect 5169 5148 5181 5151
rect 4304 5120 5181 5148
rect 4304 5108 4310 5120
rect 5169 5117 5181 5120
rect 5215 5117 5227 5151
rect 5169 5111 5227 5117
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 6564 5148 6592 5176
rect 5592 5120 6592 5148
rect 5592 5108 5598 5120
rect 6733 5015 6791 5021
rect 6733 4981 6745 5015
rect 6779 5012 6791 5015
rect 6822 5012 6828 5024
rect 6779 4984 6828 5012
rect 6779 4981 6791 4984
rect 6733 4975 6791 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 3036 4922 9844 4944
rect 3036 4870 7566 4922
rect 7618 4870 7630 4922
rect 7682 4870 7694 4922
rect 7746 4870 7758 4922
rect 7810 4870 7822 4922
rect 7874 4870 9844 4922
rect 3036 4848 9844 4870
rect 13814 4836 13820 4888
rect 13872 4876 13878 4888
rect 14090 4876 14096 4888
rect 13872 4848 14096 4876
rect 13872 4836 13878 4848
rect 14090 4836 14096 4848
rect 14148 4836 14154 4888
rect 290 4768 296 4820
rect 348 4808 354 4820
rect 2590 4808 2596 4820
rect 348 4780 2596 4808
rect 348 4768 354 4780
rect 2590 4768 2596 4780
rect 2648 4768 2654 4820
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 3970 4808 3976 4820
rect 3651 4780 3976 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 4709 4811 4767 4817
rect 4709 4777 4721 4811
rect 4755 4808 4767 4811
rect 5166 4808 5172 4820
rect 4755 4780 5172 4808
rect 4755 4777 4767 4780
rect 4709 4771 4767 4777
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5442 4808 5448 4820
rect 5307 4780 5448 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 6733 4811 6791 4817
rect 6733 4808 6745 4811
rect 6144 4780 6745 4808
rect 6144 4768 6150 4780
rect 6733 4777 6745 4780
rect 6779 4777 6791 4811
rect 7374 4808 7380 4820
rect 7335 4780 7380 4808
rect 6733 4771 6791 4777
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 8389 4811 8447 4817
rect 8389 4777 8401 4811
rect 8435 4808 8447 4811
rect 8478 4808 8484 4820
rect 8435 4780 8484 4808
rect 8435 4777 8447 4780
rect 8389 4771 8447 4777
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 9214 4808 9220 4820
rect 9175 4780 9220 4808
rect 9214 4768 9220 4780
rect 9272 4768 9278 4820
rect 750 4700 756 4752
rect 808 4740 814 4752
rect 4246 4740 4252 4752
rect 808 4712 4252 4740
rect 808 4700 814 4712
rect 4246 4700 4252 4712
rect 4304 4700 4310 4752
rect 5994 4740 6000 4752
rect 5955 4712 6000 4740
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 658 4632 664 4684
rect 716 4672 722 4684
rect 5810 4672 5816 4684
rect 716 4644 4568 4672
rect 716 4632 722 4644
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 2866 4604 2872 4616
rect 1360 4576 2872 4604
rect 1360 4564 1366 4576
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 3510 4604 3516 4616
rect 3471 4576 3516 4604
rect 3510 4564 3516 4576
rect 3568 4604 3574 4616
rect 3970 4604 3976 4616
rect 3568 4576 3976 4604
rect 3568 4564 3574 4576
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4540 4613 4568 4644
rect 5184 4644 5816 4672
rect 5184 4613 5212 4644
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 8110 4672 8116 4684
rect 7300 4644 8116 4672
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4573 5227 4607
rect 5350 4604 5356 4616
rect 5311 4576 5356 4604
rect 5169 4567 5227 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 6178 4604 6184 4616
rect 6139 4576 6184 4604
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 7300 4613 7328 4644
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 6788 4576 6837 4604
rect 6788 4564 6794 4576
rect 6825 4573 6837 4576
rect 6871 4573 6883 4607
rect 6825 4567 6883 4573
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 7432 4576 7481 4604
rect 7432 4564 7438 4576
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 8570 4604 8576 4616
rect 8531 4576 8576 4604
rect 7469 4567 7527 4573
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4604 9091 4607
rect 9398 4604 9404 4616
rect 9079 4576 9404 4604
rect 9079 4573 9091 4576
rect 9033 4567 9091 4573
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 842 4496 848 4548
rect 900 4536 906 4548
rect 2958 4536 2964 4548
rect 900 4508 2964 4536
rect 900 4496 906 4508
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 9950 4468 9956 4480
rect 8260 4440 9956 4468
rect 8260 4428 8266 4440
rect 9950 4428 9956 4440
rect 10008 4428 10014 4480
rect 3036 4378 9844 4400
rect 3036 4326 3566 4378
rect 3618 4326 3630 4378
rect 3682 4326 3694 4378
rect 3746 4326 3758 4378
rect 3810 4326 3822 4378
rect 3874 4326 8566 4378
rect 8618 4326 8630 4378
rect 8682 4326 8694 4378
rect 8746 4326 8758 4378
rect 8810 4326 8822 4378
rect 8874 4326 9844 4378
rect 3036 4304 9844 4326
rect 7009 4267 7067 4273
rect 7009 4233 7021 4267
rect 7055 4264 7067 4267
rect 7098 4264 7104 4276
rect 7055 4236 7104 4264
rect 7055 4233 7067 4236
rect 7009 4227 7067 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 7374 4224 7380 4276
rect 7432 4264 7438 4276
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 7432 4236 7573 4264
rect 7432 4224 7438 4236
rect 7561 4233 7573 4236
rect 7607 4233 7619 4267
rect 7561 4227 7619 4233
rect 3970 4156 3976 4208
rect 4028 4196 4034 4208
rect 4028 4168 4200 4196
rect 4028 4156 4034 4168
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 2832 4100 3709 4128
rect 2832 4088 2838 4100
rect 3697 4097 3709 4100
rect 3743 4097 3755 4131
rect 4062 4128 4068 4140
rect 4023 4100 4068 4128
rect 3697 4091 3755 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4172 4128 4200 4168
rect 6546 4156 6552 4208
rect 6604 4196 6610 4208
rect 7392 4196 7420 4224
rect 6604 4168 6960 4196
rect 6604 4156 6610 4168
rect 4798 4128 4804 4140
rect 4172 4100 4804 4128
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5626 4128 5632 4140
rect 4948 4100 4993 4128
rect 5587 4100 5632 4128
rect 4948 4088 4954 4100
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 6089 4131 6147 4137
rect 6089 4128 6101 4131
rect 5776 4100 6101 4128
rect 5776 4088 5782 4100
rect 6089 4097 6101 4100
rect 6135 4097 6147 4131
rect 6089 4091 6147 4097
rect 6273 4131 6331 4137
rect 6273 4097 6285 4131
rect 6319 4128 6331 4131
rect 6362 4128 6368 4140
rect 6319 4100 6368 4128
rect 6319 4097 6331 4100
rect 6273 4091 6331 4097
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6696 4100 6837 4128
rect 6696 4088 6702 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 3970 4020 3976 4072
rect 4028 4060 4034 4072
rect 4430 4060 4436 4072
rect 4028 4032 4436 4060
rect 4028 4020 4034 4032
rect 4430 4020 4436 4032
rect 4488 4020 4494 4072
rect 6932 4060 6960 4168
rect 7024 4168 7420 4196
rect 7024 4137 7052 4168
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4128 9091 4131
rect 9122 4128 9128 4140
rect 9079 4100 9128 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 7668 4060 7696 4091
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 6932 4032 7696 4060
rect 5442 3924 5448 3936
rect 5403 3896 5448 3924
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 6178 3924 6184 3936
rect 6139 3896 6184 3924
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 8202 3924 8208 3936
rect 7340 3896 8208 3924
rect 7340 3884 7346 3896
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 9214 3924 9220 3936
rect 9175 3896 9220 3924
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 3036 3834 9844 3856
rect 3036 3782 7566 3834
rect 7618 3782 7630 3834
rect 7682 3782 7694 3834
rect 7746 3782 7758 3834
rect 7810 3782 7822 3834
rect 7874 3782 9844 3834
rect 3036 3760 9844 3782
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 3605 3723 3663 3729
rect 3605 3720 3617 3723
rect 3476 3692 3617 3720
rect 3476 3680 3482 3692
rect 3605 3689 3617 3692
rect 3651 3689 3663 3723
rect 3605 3683 3663 3689
rect 4985 3723 5043 3729
rect 4985 3689 4997 3723
rect 5031 3720 5043 3723
rect 5074 3720 5080 3732
rect 5031 3692 5080 3720
rect 5031 3689 5043 3692
rect 4985 3683 5043 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 5994 3720 6000 3732
rect 5955 3692 6000 3720
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 11238 3720 11244 3732
rect 9263 3692 11244 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 4341 3655 4399 3661
rect 4341 3621 4353 3655
rect 4387 3652 4399 3655
rect 5258 3652 5264 3664
rect 4387 3624 5264 3652
rect 4387 3621 4399 3624
rect 4341 3615 4399 3621
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 6362 3544 6368 3596
rect 6420 3584 6426 3596
rect 6420 3556 7236 3584
rect 6420 3544 6426 3556
rect 2958 3476 2964 3528
rect 3016 3516 3022 3528
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 3016 3488 3525 3516
rect 3016 3476 3022 3488
rect 3513 3485 3525 3488
rect 3559 3485 3571 3519
rect 3513 3479 3571 3485
rect 3697 3519 3755 3525
rect 3697 3485 3709 3519
rect 3743 3485 3755 3519
rect 4154 3516 4160 3528
rect 4115 3488 4160 3516
rect 3697 3479 3755 3485
rect 3712 3448 3740 3479
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4798 3476 4804 3528
rect 4856 3516 4862 3528
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4856 3488 4905 3516
rect 4856 3476 4862 3488
rect 4893 3485 4905 3488
rect 4939 3516 4951 3519
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 4939 3488 6101 3516
rect 4939 3485 4951 3488
rect 4893 3479 4951 3485
rect 6089 3485 6101 3488
rect 6135 3516 6147 3519
rect 6822 3516 6828 3528
rect 6135 3488 6828 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 7006 3516 7012 3528
rect 6967 3488 7012 3516
rect 7006 3476 7012 3488
rect 7064 3476 7070 3528
rect 7208 3525 7236 3556
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 8202 3516 8208 3528
rect 8163 3488 8208 3516
rect 7193 3479 7251 3485
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 9033 3519 9091 3525
rect 9033 3516 9045 3519
rect 8996 3488 9045 3516
rect 8996 3476 9002 3488
rect 9033 3485 9045 3488
rect 9079 3485 9091 3519
rect 9033 3479 9091 3485
rect 3712 3420 4936 3448
rect 4908 3392 4936 3420
rect 4890 3340 4896 3392
rect 4948 3340 4954 3392
rect 7193 3383 7251 3389
rect 7193 3349 7205 3383
rect 7239 3380 7251 3383
rect 7926 3380 7932 3392
rect 7239 3352 7932 3380
rect 7239 3349 7251 3352
rect 7193 3343 7251 3349
rect 7926 3340 7932 3352
rect 7984 3340 7990 3392
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 8168 3352 8309 3380
rect 8168 3340 8174 3352
rect 8297 3349 8309 3352
rect 8343 3349 8355 3383
rect 8297 3343 8355 3349
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 9858 3380 9864 3392
rect 8444 3352 9864 3380
rect 8444 3340 8450 3352
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 3036 3290 9844 3312
rect 3036 3238 3566 3290
rect 3618 3238 3630 3290
rect 3682 3238 3694 3290
rect 3746 3238 3758 3290
rect 3810 3238 3822 3290
rect 3874 3238 8566 3290
rect 8618 3238 8630 3290
rect 8682 3238 8694 3290
rect 8746 3238 8758 3290
rect 8810 3238 8822 3290
rect 8874 3238 9844 3290
rect 3036 3216 9844 3238
rect 4893 3179 4951 3185
rect 4893 3145 4905 3179
rect 4939 3176 4951 3179
rect 5074 3176 5080 3188
rect 4939 3148 5080 3176
rect 4939 3145 4951 3148
rect 4893 3139 4951 3145
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 6181 3179 6239 3185
rect 6181 3145 6193 3179
rect 6227 3176 6239 3179
rect 7098 3176 7104 3188
rect 6227 3148 7104 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 7098 3136 7104 3148
rect 7156 3136 7162 3188
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 7466 3176 7472 3188
rect 7239 3148 7472 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 8018 3176 8024 3188
rect 7883 3148 8024 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 9214 3176 9220 3188
rect 9175 3148 9220 3176
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 4062 3108 4068 3120
rect 4023 3080 4068 3108
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 6914 3068 6920 3120
rect 6972 3108 6978 3120
rect 9490 3108 9496 3120
rect 6972 3080 7696 3108
rect 6972 3068 6978 3080
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 2924 3012 3617 3040
rect 2924 3000 2930 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 4706 3040 4712 3052
rect 4667 3012 4712 3040
rect 3605 3003 3663 3009
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 4890 3040 4896 3052
rect 4851 3012 4896 3040
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 5350 3040 5356 3052
rect 5311 3012 5356 3040
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3009 5595 3043
rect 5994 3040 6000 3052
rect 5955 3012 6000 3040
rect 5537 3003 5595 3009
rect 5552 2972 5580 3003
rect 5994 3000 6000 3012
rect 6052 3000 6058 3052
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 7282 3040 7288 3052
rect 7055 3012 7288 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7668 3049 7696 3080
rect 8680 3080 9496 3108
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3009 7711 3043
rect 8478 3040 8484 3052
rect 8439 3012 8484 3040
rect 7653 3003 7711 3009
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 8680 3049 8708 3080
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 9125 3043 9183 3049
rect 9125 3040 9137 3043
rect 9088 3012 9137 3040
rect 9088 3000 9094 3012
rect 9125 3009 9137 3012
rect 9171 3009 9183 3043
rect 9125 3003 9183 3009
rect 9214 3000 9220 3052
rect 9272 3040 9278 3052
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 9272 3012 9321 3040
rect 9272 3000 9278 3012
rect 9309 3009 9321 3012
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 7466 2972 7472 2984
rect 5552 2944 7472 2972
rect 7466 2932 7472 2944
rect 7524 2972 7530 2984
rect 11330 2972 11336 2984
rect 7524 2944 11336 2972
rect 7524 2932 7530 2944
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 4614 2864 4620 2916
rect 4672 2904 4678 2916
rect 4672 2876 5028 2904
rect 4672 2864 4678 2876
rect 5000 2848 5028 2876
rect 7190 2864 7196 2916
rect 7248 2904 7254 2916
rect 11238 2904 11244 2916
rect 7248 2876 11244 2904
rect 7248 2864 7254 2876
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 4982 2796 4988 2848
rect 5040 2796 5046 2848
rect 5442 2836 5448 2848
rect 5403 2808 5448 2836
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 8573 2839 8631 2845
rect 8573 2836 8585 2839
rect 8352 2808 8585 2836
rect 8352 2796 8358 2808
rect 8573 2805 8585 2808
rect 8619 2805 8631 2839
rect 8573 2799 8631 2805
rect 3036 2746 9844 2768
rect 3036 2694 7566 2746
rect 7618 2694 7630 2746
rect 7682 2694 7694 2746
rect 7746 2694 7758 2746
rect 7810 2694 7822 2746
rect 7874 2694 9844 2746
rect 3036 2672 9844 2694
rect 3142 2592 3148 2644
rect 3200 2632 3206 2644
rect 3605 2635 3663 2641
rect 3605 2632 3617 2635
rect 3200 2604 3617 2632
rect 3200 2592 3206 2604
rect 3605 2601 3617 2604
rect 3651 2601 3663 2635
rect 3605 2595 3663 2601
rect 4246 2592 4252 2644
rect 4304 2632 4310 2644
rect 4709 2635 4767 2641
rect 4709 2632 4721 2635
rect 4304 2604 4721 2632
rect 4304 2592 4310 2604
rect 4709 2601 4721 2604
rect 4755 2601 4767 2635
rect 4709 2595 4767 2601
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 9214 2632 9220 2644
rect 8619 2604 9220 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 4890 2524 4896 2576
rect 4948 2524 4954 2576
rect 5626 2524 5632 2576
rect 5684 2564 5690 2576
rect 5997 2567 6055 2573
rect 5997 2564 6009 2567
rect 5684 2536 6009 2564
rect 5684 2524 5690 2536
rect 5997 2533 6009 2536
rect 6043 2533 6055 2567
rect 5997 2527 6055 2533
rect 9125 2567 9183 2573
rect 9125 2533 9137 2567
rect 9171 2564 9183 2567
rect 9766 2564 9772 2576
rect 9171 2536 9772 2564
rect 9171 2533 9183 2536
rect 9125 2527 9183 2533
rect 9766 2524 9772 2536
rect 9824 2524 9830 2576
rect 4908 2496 4936 2524
rect 3712 2468 4936 2496
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 3712 2437 3740 2468
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 7926 2496 7932 2508
rect 5592 2468 6592 2496
rect 5592 2456 5598 2468
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 2832 2400 3525 2428
rect 2832 2388 2838 2400
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 3697 2431 3755 2437
rect 3697 2397 3709 2431
rect 3743 2397 3755 2431
rect 3697 2391 3755 2397
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2428 6147 2431
rect 6270 2428 6276 2440
rect 6135 2400 6276 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 3418 2320 3424 2372
rect 3476 2360 3482 2372
rect 4908 2360 4936 2391
rect 3476 2332 4936 2360
rect 5920 2360 5948 2391
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 6564 2437 6592 2468
rect 7208 2468 7932 2496
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 6638 2388 6644 2440
rect 6696 2428 6702 2440
rect 7208 2437 7236 2468
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 13354 2496 13360 2508
rect 8680 2468 13360 2496
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6696 2400 6745 2428
rect 6696 2388 6702 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2428 7435 2431
rect 8202 2428 8208 2440
rect 7423 2400 8208 2428
rect 7423 2397 7435 2400
rect 7377 2391 7435 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8680 2437 8708 2468
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2397 8723 2431
rect 9306 2428 9312 2440
rect 9267 2400 9312 2428
rect 8665 2391 8723 2397
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 7098 2360 7104 2372
rect 5920 2332 7104 2360
rect 3476 2320 3482 2332
rect 7098 2320 7104 2332
rect 7156 2320 7162 2372
rect 6638 2292 6644 2304
rect 6599 2264 6644 2292
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 6788 2264 7297 2292
rect 6788 2252 6794 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 3036 2202 9844 2224
rect 3036 2150 3566 2202
rect 3618 2150 3630 2202
rect 3682 2150 3694 2202
rect 3746 2150 3758 2202
rect 3810 2150 3822 2202
rect 3874 2150 8566 2202
rect 8618 2150 8630 2202
rect 8682 2150 8694 2202
rect 8746 2150 8758 2202
rect 8810 2150 8822 2202
rect 8874 2150 9844 2202
rect 3036 2128 9844 2150
rect 3697 2091 3755 2097
rect 3697 2057 3709 2091
rect 3743 2088 3755 2091
rect 3970 2088 3976 2100
rect 3743 2060 3976 2088
rect 3743 2057 3755 2060
rect 3697 2051 3755 2057
rect 3970 2048 3976 2060
rect 4028 2048 4034 2100
rect 4341 2091 4399 2097
rect 4341 2057 4353 2091
rect 4387 2088 4399 2091
rect 4982 2088 4988 2100
rect 4387 2060 4988 2088
rect 4387 2057 4399 2060
rect 4341 2051 4399 2057
rect 4982 2048 4988 2060
rect 5040 2048 5046 2100
rect 5626 2088 5632 2100
rect 5587 2060 5632 2088
rect 5626 2048 5632 2060
rect 5684 2048 5690 2100
rect 6270 2088 6276 2100
rect 6231 2060 6276 2088
rect 6270 2048 6276 2060
rect 6328 2048 6334 2100
rect 7469 2091 7527 2097
rect 7469 2057 7481 2091
rect 7515 2088 7527 2091
rect 8018 2088 8024 2100
rect 7515 2060 8024 2088
rect 7515 2057 7527 2060
rect 7469 2051 7527 2057
rect 8018 2048 8024 2060
rect 8076 2048 8082 2100
rect 8478 2048 8484 2100
rect 8536 2088 8542 2100
rect 9217 2091 9275 2097
rect 9217 2088 9229 2091
rect 8536 2060 9229 2088
rect 8536 2048 8542 2060
rect 9217 2057 9229 2060
rect 9263 2057 9275 2091
rect 9217 2051 9275 2057
rect 8110 2020 8116 2032
rect 6932 1992 8116 2020
rect 3513 1955 3571 1961
rect 3513 1921 3525 1955
rect 3559 1952 3571 1955
rect 4062 1952 4068 1964
rect 3559 1924 4068 1952
rect 3559 1921 3571 1924
rect 3513 1915 3571 1921
rect 4062 1912 4068 1924
rect 4120 1912 4126 1964
rect 4154 1912 4160 1964
rect 4212 1952 4218 1964
rect 4212 1924 4257 1952
rect 4212 1912 4218 1924
rect 4338 1912 4344 1964
rect 4396 1952 4402 1964
rect 4801 1955 4859 1961
rect 4801 1952 4813 1955
rect 4396 1924 4813 1952
rect 4396 1912 4402 1924
rect 4801 1921 4813 1924
rect 4847 1921 4859 1955
rect 4801 1915 4859 1921
rect 4890 1912 4896 1964
rect 4948 1952 4954 1964
rect 4985 1955 5043 1961
rect 4985 1952 4997 1955
rect 4948 1924 4997 1952
rect 4948 1912 4954 1924
rect 4985 1921 4997 1924
rect 5031 1921 5043 1955
rect 5442 1952 5448 1964
rect 5403 1924 5448 1952
rect 4985 1915 5043 1921
rect 5000 1884 5028 1915
rect 5442 1912 5448 1924
rect 5500 1912 5506 1964
rect 6086 1952 6092 1964
rect 6047 1924 6092 1952
rect 6086 1912 6092 1924
rect 6144 1912 6150 1964
rect 6178 1912 6184 1964
rect 6236 1952 6242 1964
rect 6273 1955 6331 1961
rect 6273 1952 6285 1955
rect 6236 1924 6285 1952
rect 6236 1912 6242 1924
rect 6273 1921 6285 1924
rect 6319 1921 6331 1955
rect 6730 1952 6736 1964
rect 6691 1924 6736 1952
rect 6273 1915 6331 1921
rect 6730 1912 6736 1924
rect 6788 1912 6794 1964
rect 6932 1961 6960 1992
rect 8110 1980 8116 1992
rect 8168 1980 8174 2032
rect 6917 1955 6975 1961
rect 6917 1921 6929 1955
rect 6963 1921 6975 1955
rect 6917 1915 6975 1921
rect 7006 1912 7012 1964
rect 7064 1952 7070 1964
rect 7377 1955 7435 1961
rect 7377 1952 7389 1955
rect 7064 1924 7389 1952
rect 7064 1912 7070 1924
rect 7377 1921 7389 1924
rect 7423 1921 7435 1955
rect 7377 1915 7435 1921
rect 9309 1955 9367 1961
rect 9309 1921 9321 1955
rect 9355 1952 9367 1955
rect 9582 1952 9588 1964
rect 9355 1924 9588 1952
rect 9355 1921 9367 1924
rect 9309 1915 9367 1921
rect 9582 1912 9588 1924
rect 9640 1912 9646 1964
rect 6196 1884 6224 1912
rect 8478 1884 8484 1896
rect 5000 1856 6224 1884
rect 8439 1856 8484 1884
rect 8478 1844 8484 1856
rect 8536 1844 8542 1896
rect 8662 1884 8668 1896
rect 8623 1856 8668 1884
rect 8662 1844 8668 1856
rect 8720 1844 8726 1896
rect 4706 1708 4712 1760
rect 4764 1748 4770 1760
rect 4893 1751 4951 1757
rect 4893 1748 4905 1751
rect 4764 1720 4905 1748
rect 4764 1708 4770 1720
rect 4893 1717 4905 1720
rect 4939 1717 4951 1751
rect 6822 1748 6828 1760
rect 6783 1720 6828 1748
rect 4893 1711 4951 1717
rect 6822 1708 6828 1720
rect 6880 1708 6886 1760
rect 3036 1658 9844 1680
rect 3036 1606 7566 1658
rect 7618 1606 7630 1658
rect 7682 1606 7694 1658
rect 7746 1606 7758 1658
rect 7810 1606 7822 1658
rect 7874 1606 9844 1658
rect 3036 1584 9844 1606
rect 106 1504 112 1556
rect 164 1544 170 1556
rect 4338 1544 4344 1556
rect 164 1516 4344 1544
rect 164 1504 170 1516
rect 4338 1504 4344 1516
rect 4396 1504 4402 1556
rect 934 1436 940 1488
rect 992 1476 998 1488
rect 2406 1476 2412 1488
rect 992 1448 2412 1476
rect 992 1436 998 1448
rect 2406 1436 2412 1448
rect 2464 1436 2470 1488
rect 1026 1368 1032 1420
rect 1084 1408 1090 1420
rect 2958 1408 2964 1420
rect 1084 1380 2964 1408
rect 1084 1368 1090 1380
rect 2958 1368 2964 1380
rect 3016 1368 3022 1420
rect 3602 1340 3608 1352
rect 3563 1312 3608 1340
rect 3602 1300 3608 1312
rect 3660 1300 3666 1352
rect 3697 1343 3755 1349
rect 3697 1309 3709 1343
rect 3743 1309 3755 1343
rect 4154 1340 4160 1352
rect 4115 1312 4160 1340
rect 3697 1303 3755 1309
rect 3234 1232 3240 1284
rect 3292 1272 3298 1284
rect 3712 1272 3740 1303
rect 4154 1300 4160 1312
rect 4212 1300 4218 1352
rect 4798 1340 4804 1352
rect 4759 1312 4804 1340
rect 4798 1300 4804 1312
rect 4856 1300 4862 1352
rect 5074 1300 5080 1352
rect 5132 1340 5138 1352
rect 5905 1343 5963 1349
rect 5905 1340 5917 1343
rect 5132 1312 5917 1340
rect 5132 1300 5138 1312
rect 5905 1309 5917 1312
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 6089 1343 6147 1349
rect 6089 1309 6101 1343
rect 6135 1340 6147 1343
rect 6178 1340 6184 1352
rect 6135 1312 6184 1340
rect 6135 1309 6147 1312
rect 6089 1303 6147 1309
rect 6178 1300 6184 1312
rect 6236 1300 6242 1352
rect 6730 1340 6736 1352
rect 6691 1312 6736 1340
rect 6730 1300 6736 1312
rect 6788 1300 6794 1352
rect 7374 1340 7380 1352
rect 7335 1312 7380 1340
rect 7374 1300 7380 1312
rect 7432 1300 7438 1352
rect 4062 1272 4068 1284
rect 3292 1244 4068 1272
rect 3292 1232 3298 1244
rect 4062 1232 4068 1244
rect 4120 1232 4126 1284
rect 6641 1275 6699 1281
rect 6641 1241 6653 1275
rect 6687 1272 6699 1275
rect 6822 1272 6828 1284
rect 6687 1244 6828 1272
rect 6687 1241 6699 1244
rect 6641 1235 6699 1241
rect 6822 1232 6828 1244
rect 6880 1232 6886 1284
rect 4338 1204 4344 1216
rect 4299 1176 4344 1204
rect 4338 1164 4344 1176
rect 4396 1164 4402 1216
rect 4890 1204 4896 1216
rect 4851 1176 4896 1204
rect 4890 1164 4896 1176
rect 4948 1164 4954 1216
rect 5902 1164 5908 1216
rect 5960 1204 5966 1216
rect 5997 1207 6055 1213
rect 5997 1204 6009 1207
rect 5960 1176 6009 1204
rect 5960 1164 5966 1176
rect 5997 1173 6009 1176
rect 6043 1173 6055 1207
rect 7282 1204 7288 1216
rect 7243 1176 7288 1204
rect 5997 1167 6055 1173
rect 7282 1164 7288 1176
rect 7340 1164 7346 1216
rect 3036 1114 9844 1136
rect 3036 1062 3566 1114
rect 3618 1062 3630 1114
rect 3682 1062 3694 1114
rect 3746 1062 3758 1114
rect 3810 1062 3822 1114
rect 3874 1062 8566 1114
rect 8618 1062 8630 1114
rect 8682 1062 8694 1114
rect 8746 1062 8758 1114
rect 8810 1062 8822 1114
rect 8874 1062 9844 1114
rect 3036 1040 9844 1062
<< via1 >>
rect 1676 15852 1728 15904
rect 2780 15852 2832 15904
rect 2566 15750 2618 15802
rect 2630 15750 2682 15802
rect 2694 15750 2746 15802
rect 2758 15750 2810 15802
rect 2822 15750 2874 15802
rect 7566 15750 7618 15802
rect 7630 15750 7682 15802
rect 7694 15750 7746 15802
rect 7758 15750 7810 15802
rect 7822 15750 7874 15802
rect 2412 15648 2464 15700
rect 6368 15648 6420 15700
rect 4712 15555 4764 15564
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 3240 15487 3292 15496
rect 3240 15453 3249 15487
rect 3249 15453 3283 15487
rect 3283 15453 3292 15487
rect 3240 15444 3292 15453
rect 2412 15376 2464 15428
rect 4068 15376 4120 15428
rect 4712 15521 4721 15555
rect 4721 15521 4755 15555
rect 4755 15521 4764 15555
rect 4712 15512 4764 15521
rect 4712 15376 4764 15428
rect 6828 15444 6880 15496
rect 8392 15487 8444 15496
rect 8392 15453 8401 15487
rect 8401 15453 8435 15487
rect 8435 15453 8444 15487
rect 8392 15444 8444 15453
rect 9036 15444 9088 15496
rect 5632 15376 5684 15428
rect 7380 15376 7432 15428
rect 8116 15419 8168 15428
rect 8116 15385 8125 15419
rect 8125 15385 8159 15419
rect 8159 15385 8168 15419
rect 8116 15376 8168 15385
rect 1308 15308 1360 15360
rect 3056 15351 3108 15360
rect 3056 15317 3065 15351
rect 3065 15317 3099 15351
rect 3099 15317 3108 15351
rect 3056 15308 3108 15317
rect 6644 15351 6696 15360
rect 6644 15317 6653 15351
rect 6653 15317 6687 15351
rect 6687 15317 6696 15351
rect 6644 15308 6696 15317
rect 9128 15351 9180 15360
rect 9128 15317 9137 15351
rect 9137 15317 9171 15351
rect 9171 15317 9180 15351
rect 9128 15308 9180 15317
rect 3566 15206 3618 15258
rect 3630 15206 3682 15258
rect 3694 15206 3746 15258
rect 3758 15206 3810 15258
rect 3822 15206 3874 15258
rect 8566 15206 8618 15258
rect 8630 15206 8682 15258
rect 8694 15206 8746 15258
rect 8758 15206 8810 15258
rect 8822 15206 8874 15258
rect 5632 15104 5684 15156
rect 1860 15036 1912 15088
rect 4160 15036 4212 15088
rect 7380 15036 7432 15088
rect 8208 15036 8260 15088
rect 2320 14968 2372 15020
rect 940 14900 992 14952
rect 3332 14968 3384 15020
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 5724 15011 5776 15020
rect 5724 14977 5733 15011
rect 5733 14977 5767 15011
rect 5767 14977 5776 15011
rect 5724 14968 5776 14977
rect 8944 15011 8996 15020
rect 8944 14977 8953 15011
rect 8953 14977 8987 15011
rect 8987 14977 8996 15011
rect 8944 14968 8996 14977
rect 1400 14832 1452 14884
rect 15936 14900 15988 14952
rect 2780 14875 2832 14884
rect 2780 14841 2789 14875
rect 2789 14841 2823 14875
rect 2823 14841 2832 14875
rect 2780 14832 2832 14841
rect 480 14764 532 14816
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 4068 14764 4120 14816
rect 4528 14764 4580 14816
rect 11428 14764 11480 14816
rect 2566 14662 2618 14714
rect 2630 14662 2682 14714
rect 2694 14662 2746 14714
rect 2758 14662 2810 14714
rect 2822 14662 2874 14714
rect 7566 14662 7618 14714
rect 7630 14662 7682 14714
rect 7694 14662 7746 14714
rect 7758 14662 7810 14714
rect 7822 14662 7874 14714
rect 13820 14696 13872 14748
rect 16212 14696 16264 14748
rect 3976 14492 4028 14544
rect 4804 14467 4856 14476
rect 4804 14433 4813 14467
rect 4813 14433 4847 14467
rect 4847 14433 4856 14467
rect 4804 14424 4856 14433
rect 5264 14467 5316 14476
rect 5264 14433 5273 14467
rect 5273 14433 5307 14467
rect 5307 14433 5316 14467
rect 5264 14424 5316 14433
rect 6460 14424 6512 14476
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 2504 14288 2556 14340
rect 4436 14331 4488 14340
rect 4436 14297 4445 14331
rect 4445 14297 4479 14331
rect 4479 14297 4488 14331
rect 4436 14288 4488 14297
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 3976 14220 4028 14272
rect 4160 14220 4212 14272
rect 5356 14288 5408 14340
rect 7380 14288 7432 14340
rect 8208 14356 8260 14408
rect 10692 14424 10744 14476
rect 16028 14424 16080 14476
rect 9496 14356 9548 14408
rect 8392 14288 8444 14340
rect 9404 14288 9456 14340
rect 10324 14288 10376 14340
rect 14096 14288 14148 14340
rect 8484 14220 8536 14272
rect 9312 14263 9364 14272
rect 9312 14229 9321 14263
rect 9321 14229 9355 14263
rect 9355 14229 9364 14263
rect 9312 14220 9364 14229
rect 3566 14118 3618 14170
rect 3630 14118 3682 14170
rect 3694 14118 3746 14170
rect 3758 14118 3810 14170
rect 3822 14118 3874 14170
rect 8566 14118 8618 14170
rect 8630 14118 8682 14170
rect 8694 14118 8746 14170
rect 8758 14118 8810 14170
rect 8822 14118 8874 14170
rect 2596 14059 2648 14068
rect 2596 14025 2605 14059
rect 2605 14025 2639 14059
rect 2639 14025 2648 14059
rect 2596 14016 2648 14025
rect 5448 14059 5500 14068
rect 5448 14025 5457 14059
rect 5457 14025 5491 14059
rect 5491 14025 5500 14059
rect 5448 14016 5500 14025
rect 9772 14016 9824 14068
rect 2780 13948 2832 14000
rect 7932 13948 7984 14000
rect 1492 13880 1544 13932
rect 2412 13880 2464 13932
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 4528 13923 4580 13932
rect 4528 13889 4537 13923
rect 4537 13889 4571 13923
rect 4571 13889 4580 13923
rect 4528 13880 4580 13889
rect 5448 13880 5500 13932
rect 7104 13923 7156 13932
rect 4896 13855 4948 13864
rect 4896 13821 4905 13855
rect 4905 13821 4939 13855
rect 4939 13821 4948 13855
rect 4896 13812 4948 13821
rect 2964 13744 3016 13796
rect 5080 13744 5132 13796
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 8484 13880 8536 13932
rect 8944 13923 8996 13932
rect 8944 13889 8953 13923
rect 8953 13889 8987 13923
rect 8987 13889 8996 13923
rect 8944 13880 8996 13889
rect 5908 13744 5960 13796
rect 2504 13676 2556 13728
rect 3056 13676 3108 13728
rect 2566 13574 2618 13626
rect 2630 13574 2682 13626
rect 2694 13574 2746 13626
rect 2758 13574 2810 13626
rect 2822 13574 2874 13626
rect 7566 13574 7618 13626
rect 7630 13574 7682 13626
rect 7694 13574 7746 13626
rect 7758 13574 7810 13626
rect 7822 13574 7874 13626
rect 5448 13336 5500 13388
rect 3056 13268 3108 13320
rect 1492 13243 1544 13252
rect 1492 13209 1501 13243
rect 1501 13209 1535 13243
rect 1535 13209 1544 13243
rect 1492 13200 1544 13209
rect 1584 13132 1636 13184
rect 5080 13268 5132 13320
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 6644 13200 6696 13252
rect 9128 13268 9180 13320
rect 12164 13200 12216 13252
rect 7288 13132 7340 13184
rect 8208 13175 8260 13184
rect 8208 13141 8217 13175
rect 8217 13141 8251 13175
rect 8251 13141 8260 13175
rect 8208 13132 8260 13141
rect 15568 13132 15620 13184
rect 3566 13030 3618 13082
rect 3630 13030 3682 13082
rect 3694 13030 3746 13082
rect 3758 13030 3810 13082
rect 3822 13030 3874 13082
rect 8566 13030 8618 13082
rect 8630 13030 8682 13082
rect 8694 13030 8746 13082
rect 8758 13030 8810 13082
rect 8822 13030 8874 13082
rect 13820 13064 13872 13116
rect 15660 13064 15712 13116
rect 8300 12971 8352 12980
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 3332 12860 3384 12912
rect 12164 12860 12216 12912
rect 16120 12860 16172 12912
rect 1400 12792 1452 12844
rect 1676 12792 1728 12844
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 4252 12792 4304 12844
rect 5264 12792 5316 12844
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 5816 12724 5868 12776
rect 6920 12724 6972 12776
rect 7288 12724 7340 12776
rect 848 12588 900 12640
rect 2964 12588 3016 12640
rect 3148 12588 3200 12640
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 15476 12792 15528 12844
rect 10140 12588 10192 12640
rect 2566 12486 2618 12538
rect 2630 12486 2682 12538
rect 2694 12486 2746 12538
rect 2758 12486 2810 12538
rect 2822 12486 2874 12538
rect 7566 12486 7618 12538
rect 7630 12486 7682 12538
rect 7694 12486 7746 12538
rect 7758 12486 7810 12538
rect 7822 12486 7874 12538
rect 13176 12520 13228 12572
rect 13912 12520 13964 12572
rect 2228 12384 2280 12436
rect 2872 12384 2924 12436
rect 6644 12384 6696 12436
rect 15016 12384 15068 12436
rect 15292 12384 15344 12436
rect 16488 12384 16540 12436
rect 10876 12316 10928 12368
rect 16396 12316 16448 12368
rect 2412 12248 2464 12300
rect 6920 12248 6972 12300
rect 8116 12248 8168 12300
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 3056 12112 3108 12164
rect 4068 12180 4120 12232
rect 4252 12180 4304 12232
rect 4712 12180 4764 12232
rect 6276 12223 6328 12232
rect 6276 12189 6285 12223
rect 6285 12189 6319 12223
rect 6319 12189 6328 12223
rect 6276 12180 6328 12189
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 4344 12112 4396 12164
rect 5908 12112 5960 12164
rect 8484 12112 8536 12164
rect 9404 12112 9456 12164
rect 1676 12044 1728 12096
rect 4068 12044 4120 12096
rect 5540 12044 5592 12096
rect 8300 12044 8352 12096
rect 9956 12044 10008 12096
rect 3566 11942 3618 11994
rect 3630 11942 3682 11994
rect 3694 11942 3746 11994
rect 3758 11942 3810 11994
rect 3822 11942 3874 11994
rect 8566 11942 8618 11994
rect 8630 11942 8682 11994
rect 8694 11942 8746 11994
rect 8758 11942 8810 11994
rect 8822 11942 8874 11994
rect 3056 11840 3108 11892
rect 8116 11883 8168 11892
rect 8116 11849 8125 11883
rect 8125 11849 8159 11883
rect 8159 11849 8168 11883
rect 8116 11840 8168 11849
rect 9036 11840 9088 11892
rect 11612 11840 11664 11892
rect 16580 11840 16632 11892
rect 3240 11772 3292 11824
rect 5816 11815 5868 11824
rect 5816 11781 5825 11815
rect 5825 11781 5859 11815
rect 5859 11781 5868 11815
rect 5816 11772 5868 11781
rect 6552 11772 6604 11824
rect 7288 11772 7340 11824
rect 8852 11815 8904 11824
rect 8852 11781 8861 11815
rect 8861 11781 8895 11815
rect 8895 11781 8904 11815
rect 8852 11772 8904 11781
rect 11428 11772 11480 11824
rect 13728 11772 13780 11824
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 8944 11704 8996 11756
rect 3240 11636 3292 11688
rect 4160 11679 4212 11688
rect 4160 11645 4169 11679
rect 4169 11645 4203 11679
rect 4203 11645 4212 11679
rect 4160 11636 4212 11645
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 15476 11568 15528 11620
rect 15752 11568 15804 11620
rect 1860 11543 1912 11552
rect 1860 11509 1869 11543
rect 1869 11509 1903 11543
rect 1903 11509 1912 11543
rect 1860 11500 1912 11509
rect 5908 11500 5960 11552
rect 7288 11500 7340 11552
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 7566 11398 7618 11450
rect 7630 11398 7682 11450
rect 7694 11398 7746 11450
rect 7758 11398 7810 11450
rect 7822 11398 7874 11450
rect 15292 11364 15344 11416
rect 16672 11364 16724 11416
rect 3332 11296 3384 11348
rect 1768 11160 1820 11212
rect 1860 11160 1912 11212
rect 4896 11203 4948 11212
rect 1860 11024 1912 11076
rect 4896 11169 4905 11203
rect 4905 11169 4939 11203
rect 4939 11169 4948 11203
rect 4896 11160 4948 11169
rect 5172 11160 5224 11212
rect 13360 11160 13412 11212
rect 15660 11228 15712 11280
rect 7104 11092 7156 11144
rect 9036 11092 9088 11144
rect 11704 11092 11756 11144
rect 13820 11092 13872 11144
rect 15476 11092 15528 11144
rect 15660 11092 15712 11144
rect 4160 11024 4212 11076
rect 5448 11024 5500 11076
rect 7196 11067 7248 11076
rect 7196 11033 7205 11067
rect 7205 11033 7239 11067
rect 7239 11033 7248 11067
rect 7196 11024 7248 11033
rect 4068 10956 4120 11008
rect 5632 10956 5684 11008
rect 8484 11024 8536 11076
rect 15476 10956 15528 11008
rect 3566 10854 3618 10906
rect 3630 10854 3682 10906
rect 3694 10854 3746 10906
rect 3758 10854 3810 10906
rect 3822 10854 3874 10906
rect 8566 10854 8618 10906
rect 8630 10854 8682 10906
rect 8694 10854 8746 10906
rect 8758 10854 8810 10906
rect 8822 10854 8874 10906
rect 15384 10888 15436 10940
rect 15936 10888 15988 10940
rect 2320 10752 2372 10804
rect 1400 10727 1452 10736
rect 1400 10693 1409 10727
rect 1409 10693 1443 10727
rect 1443 10693 1452 10727
rect 1400 10684 1452 10693
rect 4896 10752 4948 10804
rect 8024 10752 8076 10804
rect 8668 10752 8720 10804
rect 9128 10752 9180 10804
rect 15936 10752 15988 10804
rect 5724 10684 5776 10736
rect 7196 10684 7248 10736
rect 2044 10616 2096 10668
rect 2136 10616 2188 10668
rect 4620 10616 4672 10668
rect 5356 10616 5408 10668
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 6184 10616 6236 10668
rect 8300 10659 8352 10668
rect 8300 10625 8309 10659
rect 8309 10625 8343 10659
rect 8343 10625 8352 10659
rect 8300 10616 8352 10625
rect 8392 10616 8444 10668
rect 2504 10591 2556 10600
rect 2504 10557 2513 10591
rect 2513 10557 2547 10591
rect 2547 10557 2556 10591
rect 2504 10548 2556 10557
rect 7932 10548 7984 10600
rect 16304 10480 16356 10532
rect 5264 10412 5316 10464
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 6092 10412 6144 10464
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 7566 10310 7618 10362
rect 7630 10310 7682 10362
rect 7694 10310 7746 10362
rect 7758 10310 7810 10362
rect 7822 10310 7874 10362
rect 2136 10251 2188 10260
rect 2136 10217 2145 10251
rect 2145 10217 2179 10251
rect 2179 10217 2188 10251
rect 2136 10208 2188 10217
rect 8944 10251 8996 10260
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 10140 10208 10192 10260
rect 16764 10208 16816 10260
rect 1676 10072 1728 10124
rect 2228 10072 2280 10124
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 9404 10072 9456 10124
rect 3424 10004 3476 10056
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 8484 10004 8536 10056
rect 5908 9936 5960 9988
rect 6920 9936 6972 9988
rect 8208 9936 8260 9988
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 6644 9868 6696 9920
rect 6828 9868 6880 9920
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 8668 9868 8720 9920
rect 9128 9911 9180 9920
rect 9128 9877 9155 9911
rect 9155 9877 9180 9911
rect 9128 9868 9180 9877
rect 13820 9868 13872 9920
rect 15108 9868 15160 9920
rect 3566 9766 3618 9818
rect 3630 9766 3682 9818
rect 3694 9766 3746 9818
rect 3758 9766 3810 9818
rect 3822 9766 3874 9818
rect 8566 9766 8618 9818
rect 8630 9766 8682 9818
rect 8694 9766 8746 9818
rect 8758 9766 8810 9818
rect 8822 9766 8874 9818
rect 16212 9800 16264 9852
rect 11704 9732 11756 9784
rect 16856 9732 16908 9784
rect 2964 9596 3016 9648
rect 3240 9596 3292 9648
rect 4344 9596 4396 9648
rect 7380 9639 7432 9648
rect 7380 9605 7389 9639
rect 7389 9605 7423 9639
rect 7423 9605 7432 9639
rect 7380 9596 7432 9605
rect 13820 9664 13872 9716
rect 15108 9664 15160 9716
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 3976 9528 4028 9580
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 7012 9528 7064 9580
rect 15200 9528 15252 9580
rect 15476 9528 15528 9580
rect 16488 9528 16540 9580
rect 16856 9528 16908 9580
rect 2228 9460 2280 9512
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 2964 9460 3016 9512
rect 5816 9503 5868 9512
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 5816 9460 5868 9469
rect 4804 9324 4856 9376
rect 9036 9324 9088 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 7566 9222 7618 9274
rect 7630 9222 7682 9274
rect 7694 9222 7746 9274
rect 7758 9222 7810 9274
rect 7822 9222 7874 9274
rect 13820 9188 13872 9240
rect 15568 9188 15620 9240
rect 4712 9163 4764 9172
rect 4712 9129 4721 9163
rect 4721 9129 4755 9163
rect 4755 9129 4764 9163
rect 4712 9120 4764 9129
rect 1768 9027 1820 9036
rect 1768 8993 1777 9027
rect 1777 8993 1811 9027
rect 1811 8993 1820 9027
rect 1768 8984 1820 8993
rect 3056 8984 3108 9036
rect 3332 8984 3384 9036
rect 7012 8984 7064 9036
rect 1492 8959 1544 8968
rect 1492 8925 1501 8959
rect 1501 8925 1535 8959
rect 1535 8925 1544 8959
rect 1492 8916 1544 8925
rect 4160 8916 4212 8968
rect 5448 8916 5500 8968
rect 7288 8916 7340 8968
rect 9036 8959 9088 8968
rect 9036 8925 9045 8959
rect 9045 8925 9079 8959
rect 9079 8925 9088 8959
rect 9036 8916 9088 8925
rect 3332 8848 3384 8900
rect 1768 8780 1820 8832
rect 6552 8823 6604 8832
rect 6552 8789 6561 8823
rect 6561 8789 6595 8823
rect 6595 8789 6604 8823
rect 6552 8780 6604 8789
rect 9128 8823 9180 8832
rect 9128 8789 9137 8823
rect 9137 8789 9171 8823
rect 9171 8789 9180 8823
rect 9128 8780 9180 8789
rect 9588 8780 9640 8832
rect 15292 8780 15344 8832
rect 3566 8678 3618 8730
rect 3630 8678 3682 8730
rect 3694 8678 3746 8730
rect 3758 8678 3810 8730
rect 3822 8678 3874 8730
rect 8566 8678 8618 8730
rect 8630 8678 8682 8730
rect 8694 8678 8746 8730
rect 8758 8678 8810 8730
rect 8822 8678 8874 8730
rect 4804 8576 4856 8628
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 5632 8576 5684 8585
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 9496 8576 9548 8628
rect 16488 8576 16540 8628
rect 3884 8508 3936 8560
rect 9128 8551 9180 8560
rect 9128 8517 9137 8551
rect 9137 8517 9171 8551
rect 9171 8517 9180 8551
rect 9128 8508 9180 8517
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 4436 8440 4488 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 9588 8440 9640 8492
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 8208 8415 8260 8424
rect 2780 8372 2832 8381
rect 8208 8381 8217 8415
rect 8217 8381 8251 8415
rect 8251 8381 8260 8415
rect 8208 8372 8260 8381
rect 10508 8372 10560 8424
rect 15752 8372 15804 8424
rect 6460 8304 6512 8356
rect 7012 8304 7064 8356
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 7566 8134 7618 8186
rect 7630 8134 7682 8186
rect 7694 8134 7746 8186
rect 7758 8134 7810 8186
rect 7822 8134 7874 8186
rect 5264 8032 5316 8084
rect 9496 8032 9548 8084
rect 3240 7896 3292 7948
rect 1584 7828 1636 7880
rect 7380 7828 7432 7880
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 9036 7828 9088 7880
rect 3240 7803 3292 7812
rect 3240 7769 3249 7803
rect 3249 7769 3283 7803
rect 3283 7769 3292 7803
rect 3240 7760 3292 7769
rect 5264 7803 5316 7812
rect 5264 7769 5273 7803
rect 5273 7769 5307 7803
rect 5307 7769 5316 7803
rect 5264 7760 5316 7769
rect 8116 7760 8168 7812
rect 4988 7692 5040 7744
rect 7012 7692 7064 7744
rect 9128 7692 9180 7744
rect 9220 7692 9272 7744
rect 3566 7590 3618 7642
rect 3630 7590 3682 7642
rect 3694 7590 3746 7642
rect 3758 7590 3810 7642
rect 3822 7590 3874 7642
rect 8566 7590 8618 7642
rect 8630 7590 8682 7642
rect 8694 7590 8746 7642
rect 8758 7590 8810 7642
rect 8822 7590 8874 7642
rect 5356 7488 5408 7540
rect 8024 7488 8076 7540
rect 8944 7488 8996 7540
rect 1492 7420 1544 7472
rect 3424 7420 3476 7472
rect 4068 7420 4120 7472
rect 4252 7420 4304 7472
rect 4804 7420 4856 7472
rect 7104 7420 7156 7472
rect 8024 7352 8076 7404
rect 9496 7352 9548 7404
rect 3424 7284 3476 7336
rect 6368 7327 6420 7336
rect 6368 7293 6377 7327
rect 6377 7293 6411 7327
rect 6411 7293 6420 7327
rect 6368 7284 6420 7293
rect 6920 7284 6972 7336
rect 8944 7148 8996 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 7566 7046 7618 7098
rect 7630 7046 7682 7098
rect 7694 7046 7746 7098
rect 7758 7046 7810 7098
rect 7822 7046 7874 7098
rect 10784 7080 10836 7132
rect 15384 7080 15436 7132
rect 10876 6944 10928 6996
rect 16948 6944 17000 6996
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 4252 6876 4304 6928
rect 4160 6808 4212 6860
rect 4804 6808 4856 6860
rect 11152 6808 11204 6860
rect 16028 6808 16080 6860
rect 3332 6740 3384 6792
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 6092 6783 6144 6792
rect 5632 6740 5684 6749
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 7472 6740 7524 6792
rect 8116 6740 8168 6792
rect 9312 6740 9364 6792
rect 7104 6672 7156 6724
rect 8852 6672 8904 6724
rect 13176 6672 13228 6724
rect 13636 6672 13688 6724
rect 3332 6604 3384 6656
rect 5540 6604 5592 6656
rect 7932 6604 7984 6656
rect 9036 6604 9088 6656
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 3566 6502 3618 6554
rect 3630 6502 3682 6554
rect 3694 6502 3746 6554
rect 3758 6502 3810 6554
rect 3822 6502 3874 6554
rect 8566 6502 8618 6554
rect 8630 6502 8682 6554
rect 8694 6502 8746 6554
rect 8758 6502 8810 6554
rect 8822 6502 8874 6554
rect 2964 6400 3016 6452
rect 3056 6400 3108 6452
rect 3424 6400 3476 6452
rect 4160 6332 4212 6384
rect 5632 6400 5684 6452
rect 13820 6400 13872 6452
rect 15660 6400 15712 6452
rect 7380 6332 7432 6384
rect 6000 6264 6052 6316
rect 7012 6264 7064 6316
rect 9772 6264 9824 6316
rect 3332 6196 3384 6248
rect 5356 6196 5408 6248
rect 6828 6196 6880 6248
rect 13084 6196 13136 6248
rect 16856 6196 16908 6248
rect 5724 6128 5776 6180
rect 13820 6128 13872 6180
rect 15936 6128 15988 6180
rect 8852 6103 8904 6112
rect 8852 6069 8861 6103
rect 8861 6069 8895 6103
rect 8895 6069 8904 6103
rect 8852 6060 8904 6069
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 7566 5958 7618 6010
rect 7630 5958 7682 6010
rect 7694 5958 7746 6010
rect 7758 5958 7810 6010
rect 7822 5958 7874 6010
rect 2412 5856 2464 5908
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 6920 5856 6972 5908
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 2688 5788 2740 5840
rect 3424 5720 3476 5772
rect 8300 5720 8352 5772
rect 9128 5720 9180 5772
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 2320 5652 2372 5704
rect 8208 5652 8260 5704
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 3332 5584 3384 5636
rect 4160 5584 4212 5636
rect 6000 5584 6052 5636
rect 9496 5584 9548 5636
rect 13820 5584 13872 5636
rect 5540 5516 5592 5568
rect 6552 5516 6604 5568
rect 7932 5516 7984 5568
rect 8392 5516 8444 5568
rect 9036 5559 9088 5568
rect 9036 5525 9045 5559
rect 9045 5525 9079 5559
rect 9079 5525 9088 5559
rect 9036 5516 9088 5525
rect 3566 5414 3618 5466
rect 3630 5414 3682 5466
rect 3694 5414 3746 5466
rect 3758 5414 3810 5466
rect 3822 5414 3874 5466
rect 8566 5414 8618 5466
rect 8630 5414 8682 5466
rect 8694 5414 8746 5466
rect 8758 5414 8810 5466
rect 8822 5414 8874 5466
rect 112 5312 164 5364
rect 2412 5312 2464 5364
rect 4068 5355 4120 5364
rect 4068 5321 4077 5355
rect 4077 5321 4111 5355
rect 4111 5321 4120 5355
rect 4068 5312 4120 5321
rect 6460 5312 6512 5364
rect 6920 5312 6972 5364
rect 6736 5244 6788 5296
rect 9220 5287 9272 5296
rect 5264 5176 5316 5228
rect 5816 5176 5868 5228
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 9220 5253 9229 5287
rect 9229 5253 9263 5287
rect 9263 5253 9272 5287
rect 9220 5244 9272 5253
rect 6552 5176 6604 5185
rect 7932 5176 7984 5228
rect 10048 5176 10100 5228
rect 4252 5108 4304 5160
rect 5540 5108 5592 5160
rect 6828 4972 6880 5024
rect 7566 4870 7618 4922
rect 7630 4870 7682 4922
rect 7694 4870 7746 4922
rect 7758 4870 7810 4922
rect 7822 4870 7874 4922
rect 13820 4836 13872 4888
rect 14096 4836 14148 4888
rect 296 4768 348 4820
rect 2596 4768 2648 4820
rect 3976 4768 4028 4820
rect 5172 4768 5224 4820
rect 5448 4768 5500 4820
rect 6092 4768 6144 4820
rect 7380 4811 7432 4820
rect 7380 4777 7389 4811
rect 7389 4777 7423 4811
rect 7423 4777 7432 4811
rect 7380 4768 7432 4777
rect 8484 4768 8536 4820
rect 9220 4811 9272 4820
rect 9220 4777 9229 4811
rect 9229 4777 9263 4811
rect 9263 4777 9272 4811
rect 9220 4768 9272 4777
rect 756 4700 808 4752
rect 4252 4700 4304 4752
rect 6000 4743 6052 4752
rect 6000 4709 6009 4743
rect 6009 4709 6043 4743
rect 6043 4709 6052 4743
rect 6000 4700 6052 4709
rect 664 4632 716 4684
rect 1308 4564 1360 4616
rect 2872 4564 2924 4616
rect 3516 4607 3568 4616
rect 3516 4573 3525 4607
rect 3525 4573 3559 4607
rect 3559 4573 3568 4607
rect 3516 4564 3568 4573
rect 3976 4564 4028 4616
rect 5816 4632 5868 4684
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 6736 4564 6788 4616
rect 8116 4632 8168 4684
rect 7380 4564 7432 4616
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 9404 4564 9456 4616
rect 848 4496 900 4548
rect 2964 4496 3016 4548
rect 8208 4428 8260 4480
rect 9956 4428 10008 4480
rect 3566 4326 3618 4378
rect 3630 4326 3682 4378
rect 3694 4326 3746 4378
rect 3758 4326 3810 4378
rect 3822 4326 3874 4378
rect 8566 4326 8618 4378
rect 8630 4326 8682 4378
rect 8694 4326 8746 4378
rect 8758 4326 8810 4378
rect 8822 4326 8874 4378
rect 7104 4224 7156 4276
rect 7380 4224 7432 4276
rect 3976 4156 4028 4208
rect 2780 4088 2832 4140
rect 4068 4131 4120 4140
rect 4068 4097 4077 4131
rect 4077 4097 4111 4131
rect 4111 4097 4120 4131
rect 4068 4088 4120 4097
rect 6552 4156 6604 4208
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 5632 4131 5684 4140
rect 4896 4088 4948 4097
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 5724 4088 5776 4140
rect 6368 4088 6420 4140
rect 6644 4088 6696 4140
rect 3976 4020 4028 4072
rect 4436 4020 4488 4072
rect 9128 4088 9180 4140
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 7288 3884 7340 3936
rect 8208 3884 8260 3936
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 7566 3782 7618 3834
rect 7630 3782 7682 3834
rect 7694 3782 7746 3834
rect 7758 3782 7810 3834
rect 7822 3782 7874 3834
rect 3424 3680 3476 3732
rect 5080 3680 5132 3732
rect 6000 3723 6052 3732
rect 6000 3689 6009 3723
rect 6009 3689 6043 3723
rect 6043 3689 6052 3723
rect 6000 3680 6052 3689
rect 11244 3680 11296 3732
rect 5264 3612 5316 3664
rect 6368 3544 6420 3596
rect 2964 3476 3016 3528
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4804 3476 4856 3528
rect 6828 3476 6880 3528
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 8944 3476 8996 3528
rect 4896 3340 4948 3392
rect 7932 3340 7984 3392
rect 8116 3340 8168 3392
rect 8392 3340 8444 3392
rect 9864 3340 9916 3392
rect 3566 3238 3618 3290
rect 3630 3238 3682 3290
rect 3694 3238 3746 3290
rect 3758 3238 3810 3290
rect 3822 3238 3874 3290
rect 8566 3238 8618 3290
rect 8630 3238 8682 3290
rect 8694 3238 8746 3290
rect 8758 3238 8810 3290
rect 8822 3238 8874 3290
rect 5080 3136 5132 3188
rect 7104 3136 7156 3188
rect 7472 3136 7524 3188
rect 8024 3136 8076 3188
rect 9220 3179 9272 3188
rect 9220 3145 9229 3179
rect 9229 3145 9263 3179
rect 9263 3145 9272 3179
rect 9220 3136 9272 3145
rect 4068 3111 4120 3120
rect 4068 3077 4077 3111
rect 4077 3077 4111 3111
rect 4111 3077 4120 3111
rect 4068 3068 4120 3077
rect 6920 3068 6972 3120
rect 2872 3000 2924 3052
rect 4712 3043 4764 3052
rect 4712 3009 4721 3043
rect 4721 3009 4755 3043
rect 4755 3009 4764 3043
rect 4712 3000 4764 3009
rect 4896 3043 4948 3052
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 6000 3043 6052 3052
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 6000 3000 6052 3009
rect 7288 3000 7340 3052
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 9496 3068 9548 3120
rect 9036 3000 9088 3052
rect 9220 3000 9272 3052
rect 7472 2932 7524 2984
rect 11336 2932 11388 2984
rect 4620 2864 4672 2916
rect 7196 2864 7248 2916
rect 11244 2864 11296 2916
rect 4988 2796 5040 2848
rect 5448 2839 5500 2848
rect 5448 2805 5457 2839
rect 5457 2805 5491 2839
rect 5491 2805 5500 2839
rect 5448 2796 5500 2805
rect 8300 2796 8352 2848
rect 7566 2694 7618 2746
rect 7630 2694 7682 2746
rect 7694 2694 7746 2746
rect 7758 2694 7810 2746
rect 7822 2694 7874 2746
rect 3148 2592 3200 2644
rect 4252 2592 4304 2644
rect 9220 2592 9272 2644
rect 4896 2524 4948 2576
rect 5632 2524 5684 2576
rect 9772 2524 9824 2576
rect 2780 2388 2832 2440
rect 5540 2456 5592 2508
rect 3424 2320 3476 2372
rect 6276 2388 6328 2440
rect 6644 2388 6696 2440
rect 7932 2456 7984 2508
rect 8208 2388 8260 2440
rect 13360 2456 13412 2508
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 7104 2320 7156 2372
rect 6644 2295 6696 2304
rect 6644 2261 6653 2295
rect 6653 2261 6687 2295
rect 6687 2261 6696 2295
rect 6644 2252 6696 2261
rect 6736 2252 6788 2304
rect 3566 2150 3618 2202
rect 3630 2150 3682 2202
rect 3694 2150 3746 2202
rect 3758 2150 3810 2202
rect 3822 2150 3874 2202
rect 8566 2150 8618 2202
rect 8630 2150 8682 2202
rect 8694 2150 8746 2202
rect 8758 2150 8810 2202
rect 8822 2150 8874 2202
rect 3976 2048 4028 2100
rect 4988 2048 5040 2100
rect 5632 2091 5684 2100
rect 5632 2057 5641 2091
rect 5641 2057 5675 2091
rect 5675 2057 5684 2091
rect 5632 2048 5684 2057
rect 6276 2091 6328 2100
rect 6276 2057 6285 2091
rect 6285 2057 6319 2091
rect 6319 2057 6328 2091
rect 6276 2048 6328 2057
rect 8024 2048 8076 2100
rect 8484 2048 8536 2100
rect 4068 1912 4120 1964
rect 4160 1955 4212 1964
rect 4160 1921 4169 1955
rect 4169 1921 4203 1955
rect 4203 1921 4212 1955
rect 4160 1912 4212 1921
rect 4344 1912 4396 1964
rect 4896 1912 4948 1964
rect 5448 1955 5500 1964
rect 5448 1921 5457 1955
rect 5457 1921 5491 1955
rect 5491 1921 5500 1955
rect 5448 1912 5500 1921
rect 6092 1955 6144 1964
rect 6092 1921 6101 1955
rect 6101 1921 6135 1955
rect 6135 1921 6144 1955
rect 6092 1912 6144 1921
rect 6184 1912 6236 1964
rect 6736 1955 6788 1964
rect 6736 1921 6745 1955
rect 6745 1921 6779 1955
rect 6779 1921 6788 1955
rect 6736 1912 6788 1921
rect 8116 1980 8168 2032
rect 7012 1912 7064 1964
rect 9588 1912 9640 1964
rect 8484 1887 8536 1896
rect 8484 1853 8493 1887
rect 8493 1853 8527 1887
rect 8527 1853 8536 1887
rect 8484 1844 8536 1853
rect 8668 1887 8720 1896
rect 8668 1853 8677 1887
rect 8677 1853 8711 1887
rect 8711 1853 8720 1887
rect 8668 1844 8720 1853
rect 4712 1708 4764 1760
rect 6828 1751 6880 1760
rect 6828 1717 6837 1751
rect 6837 1717 6871 1751
rect 6871 1717 6880 1751
rect 6828 1708 6880 1717
rect 7566 1606 7618 1658
rect 7630 1606 7682 1658
rect 7694 1606 7746 1658
rect 7758 1606 7810 1658
rect 7822 1606 7874 1658
rect 112 1504 164 1556
rect 4344 1504 4396 1556
rect 940 1436 992 1488
rect 2412 1436 2464 1488
rect 1032 1368 1084 1420
rect 2964 1368 3016 1420
rect 3608 1343 3660 1352
rect 3608 1309 3617 1343
rect 3617 1309 3651 1343
rect 3651 1309 3660 1343
rect 3608 1300 3660 1309
rect 4160 1343 4212 1352
rect 3240 1232 3292 1284
rect 4160 1309 4169 1343
rect 4169 1309 4203 1343
rect 4203 1309 4212 1343
rect 4160 1300 4212 1309
rect 4804 1343 4856 1352
rect 4804 1309 4813 1343
rect 4813 1309 4847 1343
rect 4847 1309 4856 1343
rect 4804 1300 4856 1309
rect 5080 1300 5132 1352
rect 6184 1300 6236 1352
rect 6736 1343 6788 1352
rect 6736 1309 6745 1343
rect 6745 1309 6779 1343
rect 6779 1309 6788 1343
rect 6736 1300 6788 1309
rect 7380 1343 7432 1352
rect 7380 1309 7389 1343
rect 7389 1309 7423 1343
rect 7423 1309 7432 1343
rect 7380 1300 7432 1309
rect 4068 1232 4120 1284
rect 6828 1232 6880 1284
rect 4344 1207 4396 1216
rect 4344 1173 4353 1207
rect 4353 1173 4387 1207
rect 4387 1173 4396 1207
rect 4344 1164 4396 1173
rect 4896 1207 4948 1216
rect 4896 1173 4905 1207
rect 4905 1173 4939 1207
rect 4939 1173 4948 1207
rect 4896 1164 4948 1173
rect 5908 1164 5960 1216
rect 7288 1207 7340 1216
rect 7288 1173 7297 1207
rect 7297 1173 7331 1207
rect 7331 1173 7340 1207
rect 7288 1164 7340 1173
rect 3566 1062 3618 1114
rect 3630 1062 3682 1114
rect 3694 1062 3746 1114
rect 3758 1062 3810 1114
rect 3822 1062 3874 1114
rect 8566 1062 8618 1114
rect 8630 1062 8682 1114
rect 8694 1062 8746 1114
rect 8758 1062 8810 1114
rect 8822 1062 8874 1114
<< metal2 >>
rect 938 16200 994 17000
rect 1398 16200 1454 17000
rect 1858 16200 1914 17000
rect 2318 16200 2374 17000
rect 2410 16960 2466 16969
rect 2410 16895 2466 16904
rect 952 14958 980 16200
rect 1214 15600 1270 15609
rect 1214 15535 1270 15544
rect 940 14952 992 14958
rect 110 14920 166 14929
rect 940 14894 992 14900
rect 110 14855 166 14864
rect 18 12880 74 12889
rect 18 12815 74 12824
rect 32 5681 60 12815
rect 18 5672 74 5681
rect 18 5607 74 5616
rect 124 5370 152 14855
rect 480 14816 532 14822
rect 480 14758 532 14764
rect 386 14104 442 14113
rect 386 14039 442 14048
rect 294 13832 350 13841
rect 294 13767 350 13776
rect 202 11112 258 11121
rect 202 11047 258 11056
rect 112 5364 164 5370
rect 112 5306 164 5312
rect 110 1592 166 1601
rect 110 1527 112 1536
rect 164 1527 166 1536
rect 112 1498 164 1504
rect 216 1465 244 11047
rect 308 4826 336 13767
rect 296 4820 348 4826
rect 296 4762 348 4768
rect 202 1456 258 1465
rect 202 1391 258 1400
rect 400 921 428 14039
rect 492 1601 520 14758
rect 662 14512 718 14521
rect 662 14447 718 14456
rect 570 14376 626 14385
rect 570 14311 626 14320
rect 478 1592 534 1601
rect 478 1527 534 1536
rect 584 1193 612 14311
rect 676 4690 704 14447
rect 754 13288 810 13297
rect 754 13223 810 13232
rect 768 4758 796 13223
rect 848 12640 900 12646
rect 848 12582 900 12588
rect 756 4752 808 4758
rect 756 4694 808 4700
rect 664 4684 716 4690
rect 664 4626 716 4632
rect 860 4554 888 12582
rect 938 12472 994 12481
rect 1228 12434 1256 15535
rect 1308 15360 1360 15366
rect 1308 15302 1360 15308
rect 938 12407 994 12416
rect 848 4548 900 4554
rect 848 4490 900 4496
rect 952 1494 980 12407
rect 1044 12406 1256 12434
rect 940 1488 992 1494
rect 940 1430 992 1436
rect 1044 1426 1072 12406
rect 1122 8392 1178 8401
rect 1122 8327 1178 8336
rect 1032 1420 1084 1426
rect 1032 1362 1084 1368
rect 1136 1329 1164 8327
rect 1320 4622 1348 15302
rect 1412 14890 1440 16200
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1400 14884 1452 14890
rect 1400 14826 1452 14832
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 13938 1532 14214
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1492 13252 1544 13258
rect 1492 13194 1544 13200
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 10742 1440 12786
rect 1504 11665 1532 13194
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 12481 1624 13126
rect 1688 12850 1716 15846
rect 1768 15496 1820 15502
rect 1766 15464 1768 15473
rect 1820 15464 1822 15473
rect 1766 15399 1822 15408
rect 1872 15094 1900 16200
rect 2332 15178 2360 16200
rect 2424 15706 2452 16895
rect 2778 16200 2834 17000
rect 3238 16200 3294 17000
rect 3436 16238 3648 16266
rect 2792 15910 2820 16200
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2566 15804 2874 15813
rect 2566 15802 2572 15804
rect 2628 15802 2652 15804
rect 2708 15802 2732 15804
rect 2788 15802 2812 15804
rect 2868 15802 2874 15804
rect 2628 15750 2630 15802
rect 2810 15750 2812 15802
rect 2566 15748 2572 15750
rect 2628 15748 2652 15750
rect 2708 15748 2732 15750
rect 2788 15748 2812 15750
rect 2868 15748 2874 15750
rect 2566 15739 2874 15748
rect 2412 15700 2464 15706
rect 3252 15688 3280 16200
rect 2412 15642 2464 15648
rect 3160 15660 3280 15688
rect 2412 15428 2464 15434
rect 2412 15370 2464 15376
rect 2240 15150 2360 15178
rect 1860 15088 1912 15094
rect 1860 15030 1912 15036
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1582 12472 1638 12481
rect 1872 12458 1900 15030
rect 1582 12407 1638 12416
rect 1780 12430 1900 12458
rect 2240 12442 2268 15150
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2228 12436 2280 12442
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1490 11656 1546 11665
rect 1490 11591 1546 11600
rect 1504 11098 1532 11591
rect 1504 11070 1624 11098
rect 1400 10736 1452 10742
rect 1400 10678 1452 10684
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1504 7478 1532 8910
rect 1596 7886 1624 11070
rect 1688 10130 1716 12038
rect 1780 11218 1808 12430
rect 2228 12378 2280 12384
rect 2332 12322 2360 14962
rect 2424 14498 2452 15370
rect 3056 15360 3108 15366
rect 3054 15328 3056 15337
rect 3108 15328 3110 15337
rect 3054 15263 3110 15272
rect 2778 14920 2834 14929
rect 2778 14855 2780 14864
rect 2832 14855 2834 14864
rect 2780 14826 2832 14832
rect 2566 14716 2874 14725
rect 2566 14714 2572 14716
rect 2628 14714 2652 14716
rect 2708 14714 2732 14716
rect 2788 14714 2812 14716
rect 2868 14714 2874 14716
rect 2628 14662 2630 14714
rect 2810 14662 2812 14714
rect 2566 14660 2572 14662
rect 2628 14660 2652 14662
rect 2708 14660 2732 14662
rect 2788 14660 2812 14662
rect 2868 14660 2874 14662
rect 2566 14651 2874 14660
rect 2424 14470 2636 14498
rect 2504 14340 2556 14346
rect 2504 14282 2556 14288
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2240 12294 2360 12322
rect 2424 12306 2452 13874
rect 2516 13734 2544 14282
rect 2608 14074 2636 14470
rect 2778 14104 2834 14113
rect 2596 14068 2648 14074
rect 2778 14039 2834 14048
rect 2596 14010 2648 14016
rect 2608 13977 2636 14010
rect 2792 14006 2820 14039
rect 2780 14000 2832 14006
rect 2594 13968 2650 13977
rect 2780 13942 2832 13948
rect 2594 13903 2650 13912
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3068 13841 3096 13874
rect 3054 13832 3110 13841
rect 2964 13796 3016 13802
rect 3054 13767 3110 13776
rect 2964 13738 3016 13744
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2566 13628 2874 13637
rect 2566 13626 2572 13628
rect 2628 13626 2652 13628
rect 2708 13626 2732 13628
rect 2788 13626 2812 13628
rect 2868 13626 2874 13628
rect 2628 13574 2630 13626
rect 2810 13574 2812 13626
rect 2566 13572 2572 13574
rect 2628 13572 2652 13574
rect 2708 13572 2732 13574
rect 2788 13572 2812 13574
rect 2868 13572 2874 13574
rect 2566 13563 2874 13572
rect 2976 12850 3004 13738
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 3068 13326 3096 13670
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2596 12776 2648 12782
rect 2594 12744 2596 12753
rect 2648 12744 2650 12753
rect 2594 12679 2650 12688
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2566 12540 2874 12549
rect 2566 12538 2572 12540
rect 2628 12538 2652 12540
rect 2708 12538 2732 12540
rect 2788 12538 2812 12540
rect 2868 12538 2874 12540
rect 2628 12486 2630 12538
rect 2810 12486 2812 12538
rect 2566 12484 2572 12486
rect 2628 12484 2652 12486
rect 2708 12484 2732 12486
rect 2788 12484 2812 12486
rect 2868 12484 2874 12486
rect 2566 12475 2874 12484
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2412 12300 2464 12306
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11218 1900 11494
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1688 9058 1716 10066
rect 1688 9042 1808 9058
rect 1688 9036 1820 9042
rect 1688 9030 1768 9036
rect 1768 8978 1820 8984
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8498 1808 8774
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1492 7472 1544 7478
rect 1492 7414 1544 7420
rect 1504 6866 1532 7414
rect 1780 6866 1808 8434
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1308 4616 1360 4622
rect 1872 4593 1900 11018
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2056 10169 2084 10610
rect 2148 10266 2176 10610
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2042 10160 2098 10169
rect 2240 10130 2268 12294
rect 2412 12242 2464 12248
rect 2884 11642 2912 12378
rect 2976 11778 3004 12582
rect 3068 12170 3096 13262
rect 3160 12646 3188 15660
rect 3238 15600 3294 15609
rect 3238 15535 3294 15544
rect 3252 15502 3280 15535
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3252 12238 3280 14350
rect 3344 13716 3372 14962
rect 3436 14056 3464 16238
rect 3620 16130 3648 16238
rect 3698 16200 3754 17000
rect 4066 16688 4122 16697
rect 4066 16623 4122 16632
rect 3712 16130 3740 16200
rect 3620 16102 3740 16130
rect 4080 15434 4108 16623
rect 4158 16200 4214 17000
rect 4618 16200 4674 17000
rect 5078 16200 5134 17000
rect 5538 16200 5594 17000
rect 5998 16200 6054 17000
rect 6366 16824 6422 16833
rect 6366 16759 6422 16768
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4066 15328 4122 15337
rect 3566 15260 3874 15269
rect 4066 15263 4122 15272
rect 3566 15258 3572 15260
rect 3628 15258 3652 15260
rect 3708 15258 3732 15260
rect 3788 15258 3812 15260
rect 3868 15258 3874 15260
rect 3628 15206 3630 15258
rect 3810 15206 3812 15258
rect 3566 15204 3572 15206
rect 3628 15204 3652 15206
rect 3708 15204 3732 15206
rect 3788 15204 3812 15206
rect 3868 15204 3874 15206
rect 3566 15195 3874 15204
rect 4080 15026 4108 15263
rect 4172 15178 4200 16200
rect 4172 15150 4384 15178
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 4068 15020 4120 15026
rect 3988 14980 4068 15008
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14385 3648 14758
rect 3988 14550 4016 14980
rect 4068 14962 4120 14968
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 3606 14376 3662 14385
rect 3606 14311 3662 14320
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 3566 14172 3874 14181
rect 3566 14170 3572 14172
rect 3628 14170 3652 14172
rect 3708 14170 3732 14172
rect 3788 14170 3812 14172
rect 3868 14170 3874 14172
rect 3628 14118 3630 14170
rect 3810 14118 3812 14170
rect 3566 14116 3572 14118
rect 3628 14116 3652 14118
rect 3708 14116 3732 14118
rect 3788 14116 3812 14118
rect 3868 14116 3874 14118
rect 3566 14107 3874 14116
rect 3436 14028 3556 14056
rect 3344 13688 3464 13716
rect 3332 12912 3384 12918
rect 3330 12880 3332 12889
rect 3384 12880 3386 12889
rect 3330 12815 3386 12824
rect 3330 12608 3386 12617
rect 3330 12543 3386 12552
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 3068 11898 3096 12106
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 3252 11830 3280 12174
rect 3240 11824 3292 11830
rect 2976 11750 3096 11778
rect 3240 11766 3292 11772
rect 2884 11614 3004 11642
rect 2566 11452 2874 11461
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11387 2874 11396
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2042 10095 2098 10104
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 2332 9738 2360 10746
rect 2504 10600 2556 10606
rect 2502 10568 2504 10577
rect 2556 10568 2558 10577
rect 2502 10503 2558 10512
rect 2566 10364 2874 10373
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10299 2874 10308
rect 2148 9710 2360 9738
rect 1950 5808 2006 5817
rect 1950 5743 2006 5752
rect 1964 5710 1992 5743
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 2148 5409 2176 9710
rect 2976 9654 3004 11614
rect 3068 10305 3096 11750
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3054 10296 3110 10305
rect 3054 10231 3110 10240
rect 3146 10024 3202 10033
rect 3252 10010 3280 11630
rect 3344 11354 3372 12543
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3436 11257 3464 13688
rect 3528 13433 3556 14028
rect 3514 13424 3570 13433
rect 3514 13359 3570 13368
rect 3566 13084 3874 13093
rect 3566 13082 3572 13084
rect 3628 13082 3652 13084
rect 3708 13082 3732 13084
rect 3788 13082 3812 13084
rect 3868 13082 3874 13084
rect 3628 13030 3630 13082
rect 3810 13030 3812 13082
rect 3566 13028 3572 13030
rect 3628 13028 3652 13030
rect 3708 13028 3732 13030
rect 3788 13028 3812 13030
rect 3868 13028 3874 13030
rect 3566 13019 3874 13028
rect 3566 11996 3874 12005
rect 3566 11994 3572 11996
rect 3628 11994 3652 11996
rect 3708 11994 3732 11996
rect 3788 11994 3812 11996
rect 3868 11994 3874 11996
rect 3628 11942 3630 11994
rect 3810 11942 3812 11994
rect 3566 11940 3572 11942
rect 3628 11940 3652 11942
rect 3708 11940 3732 11942
rect 3788 11940 3812 11942
rect 3868 11940 3874 11942
rect 3566 11931 3874 11940
rect 3422 11248 3478 11257
rect 3422 11183 3478 11192
rect 3566 10908 3874 10917
rect 3566 10906 3572 10908
rect 3628 10906 3652 10908
rect 3708 10906 3732 10908
rect 3788 10906 3812 10908
rect 3868 10906 3874 10908
rect 3628 10854 3630 10906
rect 3810 10854 3812 10906
rect 3566 10852 3572 10854
rect 3628 10852 3652 10854
rect 3708 10852 3732 10854
rect 3788 10852 3812 10854
rect 3868 10852 3874 10854
rect 3566 10843 3874 10852
rect 3424 10056 3476 10062
rect 3252 9982 3372 10010
rect 3424 9998 3476 10004
rect 3146 9959 3202 9968
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2228 9512 2280 9518
rect 2688 9512 2740 9518
rect 2228 9454 2280 9460
rect 2686 9480 2688 9489
rect 2964 9512 3016 9518
rect 2740 9480 2742 9489
rect 2134 5400 2190 5409
rect 2134 5335 2190 5344
rect 1308 4558 1360 4564
rect 1858 4584 1914 4593
rect 1858 4519 1914 4528
rect 2240 4536 2268 9454
rect 2964 9454 3016 9460
rect 2686 9415 2742 9424
rect 2566 9276 2874 9285
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9211 2874 9220
rect 2780 8424 2832 8430
rect 2778 8392 2780 8401
rect 2832 8392 2834 8401
rect 2778 8327 2834 8336
rect 2566 8188 2874 8197
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8123 2874 8132
rect 2318 7848 2374 7857
rect 2318 7783 2374 7792
rect 2332 5710 2360 7783
rect 2566 7100 2874 7109
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7035 2874 7044
rect 2976 6458 3004 9454
rect 3068 9217 3096 9522
rect 3054 9208 3110 9217
rect 3054 9143 3110 9152
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 3068 6458 3096 8978
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2410 6352 2466 6361
rect 2410 6287 2466 6296
rect 2424 5914 2452 6287
rect 3054 6080 3110 6089
rect 2566 6012 2874 6021
rect 3054 6015 3110 6024
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5947 2874 5956
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2502 5672 2558 5681
rect 2502 5607 2558 5616
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2240 4508 2360 4536
rect 2332 4026 2360 4508
rect 2424 4185 2452 5306
rect 2410 4176 2466 4185
rect 2410 4111 2466 4120
rect 2410 4040 2466 4049
rect 2332 3998 2410 4026
rect 2410 3975 2466 3984
rect 2516 3890 2544 5607
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2424 3862 2544 3890
rect 2424 2774 2452 3862
rect 2608 3777 2636 4762
rect 2700 4162 2728 5782
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2700 4146 2820 4162
rect 2700 4140 2832 4146
rect 2700 4134 2780 4140
rect 2780 4082 2832 4088
rect 2686 4040 2742 4049
rect 2686 3975 2742 3984
rect 2594 3768 2650 3777
rect 2594 3703 2650 3712
rect 2700 3641 2728 3975
rect 2686 3632 2742 3641
rect 2686 3567 2742 3576
rect 2884 3058 2912 4558
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2976 3534 3004 4490
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2332 2746 2452 2774
rect 3068 2774 3096 6015
rect 3160 3097 3188 9959
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3252 9761 3280 9862
rect 3238 9752 3294 9761
rect 3238 9687 3294 9696
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3252 8265 3280 9590
rect 3344 9042 3372 9982
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3238 8256 3294 8265
rect 3238 8191 3294 8200
rect 3252 7954 3280 8191
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3252 7313 3280 7754
rect 3238 7304 3294 7313
rect 3238 7239 3294 7248
rect 3146 3088 3202 3097
rect 3146 3023 3202 3032
rect 3068 2746 3188 2774
rect 2332 2530 2360 2746
rect 3160 2650 3188 2746
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 2410 2544 2466 2553
rect 2332 2502 2410 2530
rect 2410 2479 2466 2488
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2410 1728 2466 1737
rect 2410 1663 2466 1672
rect 1858 1592 1914 1601
rect 2318 1592 2374 1601
rect 1914 1550 2318 1578
rect 1858 1527 1914 1536
rect 2318 1527 2374 1536
rect 2424 1494 2452 1663
rect 2412 1488 2464 1494
rect 2792 1465 2820 2382
rect 2412 1430 2464 1436
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 2962 1456 3018 1465
rect 2962 1391 2964 1400
rect 3016 1391 3018 1400
rect 2964 1362 3016 1368
rect 1122 1320 1178 1329
rect 3252 1290 3280 7239
rect 3344 6798 3372 8842
rect 3436 7478 3464 9998
rect 3566 9820 3874 9829
rect 3566 9818 3572 9820
rect 3628 9818 3652 9820
rect 3708 9818 3732 9820
rect 3788 9818 3812 9820
rect 3868 9818 3874 9820
rect 3628 9766 3630 9818
rect 3810 9766 3812 9818
rect 3566 9764 3572 9766
rect 3628 9764 3652 9766
rect 3708 9764 3732 9766
rect 3788 9764 3812 9766
rect 3868 9764 3874 9766
rect 3566 9755 3874 9764
rect 3988 9586 4016 14214
rect 4080 12238 4108 14758
rect 4172 14278 4200 15030
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4250 13288 4306 13297
rect 4250 13223 4306 13232
rect 4264 12850 4292 13223
rect 4356 12889 4384 15150
rect 4632 14906 4660 16200
rect 4710 15600 4766 15609
rect 4710 15535 4712 15544
rect 4764 15535 4766 15544
rect 4712 15506 4764 15512
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4448 14878 4660 14906
rect 4448 14346 4476 14878
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 4342 12880 4398 12889
rect 4252 12844 4304 12850
rect 4342 12815 4398 12824
rect 4252 12786 4304 12792
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4068 12096 4120 12102
rect 4066 12064 4068 12073
rect 4120 12064 4122 12073
rect 4066 11999 4122 12008
rect 4160 11688 4212 11694
rect 4158 11656 4160 11665
rect 4212 11656 4214 11665
rect 4158 11591 4214 11600
rect 4158 11112 4214 11121
rect 4158 11047 4160 11056
rect 4212 11047 4214 11056
rect 4160 11018 4212 11024
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10130 4108 10950
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4264 9738 4292 12174
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 4080 9710 4292 9738
rect 4356 9738 4384 12106
rect 4448 10033 4476 14282
rect 4540 13938 4568 14758
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4724 12322 4752 15370
rect 4802 14512 4858 14521
rect 4802 14447 4804 14456
rect 4856 14447 4858 14456
rect 4804 14418 4856 14424
rect 4896 13864 4948 13870
rect 4894 13832 4896 13841
rect 4948 13832 4950 13841
rect 5092 13802 5120 16200
rect 5552 16130 5580 16200
rect 5552 16102 5764 16130
rect 5262 15464 5318 15473
rect 5262 15399 5318 15408
rect 5632 15428 5684 15434
rect 5276 14482 5304 15399
rect 5632 15370 5684 15376
rect 5644 15162 5672 15370
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5736 15026 5764 16102
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5446 14512 5502 14521
rect 5264 14476 5316 14482
rect 5446 14447 5502 14456
rect 5264 14418 5316 14424
rect 4894 13767 4950 13776
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 12434 4936 12582
rect 4908 12406 5028 12434
rect 4894 12336 4950 12345
rect 4724 12294 4844 12322
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4434 10024 4490 10033
rect 4434 9959 4490 9968
rect 4356 9710 4476 9738
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3566 8732 3874 8741
rect 3566 8730 3572 8732
rect 3628 8730 3652 8732
rect 3708 8730 3732 8732
rect 3788 8730 3812 8732
rect 3868 8730 3874 8732
rect 3628 8678 3630 8730
rect 3810 8678 3812 8730
rect 3566 8676 3572 8678
rect 3628 8676 3652 8678
rect 3708 8676 3732 8678
rect 3788 8676 3812 8678
rect 3868 8676 3874 8678
rect 3566 8667 3874 8676
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3896 8401 3924 8502
rect 3882 8392 3938 8401
rect 3882 8327 3938 8336
rect 4080 7698 4108 9710
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 3988 7670 4108 7698
rect 3566 7644 3874 7653
rect 3566 7642 3572 7644
rect 3628 7642 3652 7644
rect 3708 7642 3732 7644
rect 3788 7642 3812 7644
rect 3868 7642 3874 7644
rect 3628 7590 3630 7642
rect 3810 7590 3812 7642
rect 3566 7588 3572 7590
rect 3628 7588 3652 7590
rect 3708 7588 3732 7590
rect 3788 7588 3812 7590
rect 3868 7588 3874 7590
rect 3566 7579 3874 7588
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3436 7342 3464 7414
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3344 6254 3372 6598
rect 3436 6458 3464 7278
rect 3566 6556 3874 6565
rect 3566 6554 3572 6556
rect 3628 6554 3652 6556
rect 3708 6554 3732 6556
rect 3788 6554 3812 6556
rect 3868 6554 3874 6556
rect 3628 6502 3630 6554
rect 3810 6502 3812 6554
rect 3566 6500 3572 6502
rect 3628 6500 3652 6502
rect 3708 6500 3732 6502
rect 3788 6500 3812 6502
rect 3868 6500 3874 6502
rect 3566 6491 3874 6500
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3344 5642 3372 6190
rect 3436 5778 3464 6394
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3422 5672 3478 5681
rect 3332 5636 3384 5642
rect 3422 5607 3478 5616
rect 3332 5578 3384 5584
rect 3330 5400 3386 5409
rect 3330 5335 3386 5344
rect 3344 3913 3372 5335
rect 3330 3904 3386 3913
rect 3330 3839 3386 3848
rect 3436 3738 3464 5607
rect 3566 5468 3874 5477
rect 3566 5466 3572 5468
rect 3628 5466 3652 5468
rect 3708 5466 3732 5468
rect 3788 5466 3812 5468
rect 3868 5466 3874 5468
rect 3628 5414 3630 5466
rect 3810 5414 3812 5466
rect 3566 5412 3572 5414
rect 3628 5412 3652 5414
rect 3708 5412 3732 5414
rect 3788 5412 3812 5414
rect 3868 5412 3874 5414
rect 3566 5403 3874 5412
rect 3988 4826 4016 7670
rect 4172 7562 4200 8910
rect 4080 7534 4200 7562
rect 4080 7478 4108 7534
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4066 7032 4122 7041
rect 4066 6967 4122 6976
rect 4080 5370 4108 6967
rect 4264 6934 4292 7414
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4172 6390 4200 6802
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 4172 5642 4200 6326
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4264 5166 4292 6870
rect 4356 5681 4384 9590
rect 4448 9353 4476 9710
rect 4434 9344 4490 9353
rect 4434 9279 4490 9288
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4342 5672 4398 5681
rect 4342 5607 4398 5616
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 4252 4752 4304 4758
rect 3514 4720 3570 4729
rect 4252 4694 4304 4700
rect 3514 4655 3570 4664
rect 3528 4622 3556 4655
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3566 4380 3874 4389
rect 3566 4378 3572 4380
rect 3628 4378 3652 4380
rect 3708 4378 3732 4380
rect 3788 4378 3812 4380
rect 3868 4378 3874 4380
rect 3628 4326 3630 4378
rect 3810 4326 3812 4378
rect 3566 4324 3572 4326
rect 3628 4324 3652 4326
rect 3708 4324 3732 4326
rect 3788 4324 3812 4326
rect 3868 4324 3874 4326
rect 3566 4315 3874 4324
rect 3988 4214 4016 4558
rect 4158 4448 4214 4457
rect 4158 4383 4214 4392
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 4066 4176 4122 4185
rect 4066 4111 4068 4120
rect 4120 4111 4122 4120
rect 4068 4082 4120 4088
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 4066 4040 4122 4049
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3566 3292 3874 3301
rect 3566 3290 3572 3292
rect 3628 3290 3652 3292
rect 3708 3290 3732 3292
rect 3788 3290 3812 3292
rect 3868 3290 3874 3292
rect 3628 3238 3630 3290
rect 3810 3238 3812 3290
rect 3566 3236 3572 3238
rect 3628 3236 3652 3238
rect 3708 3236 3732 3238
rect 3788 3236 3812 3238
rect 3868 3236 3874 3238
rect 3566 3227 3874 3236
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 1122 1255 1178 1264
rect 3240 1284 3292 1290
rect 3240 1226 3292 1232
rect 3436 1193 3464 2314
rect 3566 2204 3874 2213
rect 3566 2202 3572 2204
rect 3628 2202 3652 2204
rect 3708 2202 3732 2204
rect 3788 2202 3812 2204
rect 3868 2202 3874 2204
rect 3628 2150 3630 2202
rect 3810 2150 3812 2202
rect 3566 2148 3572 2150
rect 3628 2148 3652 2150
rect 3708 2148 3732 2150
rect 3788 2148 3812 2150
rect 3868 2148 3874 2150
rect 3566 2139 3874 2148
rect 3988 2106 4016 4014
rect 4066 3975 4122 3984
rect 4080 3126 4108 3975
rect 4172 3534 4200 4383
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4066 2680 4122 2689
rect 4264 2650 4292 4694
rect 4448 4078 4476 8434
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4632 2922 4660 10610
rect 4724 9178 4752 12174
rect 4816 9382 4844 12294
rect 4894 12271 4950 12280
rect 4908 11218 4936 12271
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 5000 11121 5028 12406
rect 4986 11112 5042 11121
rect 4986 11047 5042 11056
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4908 10713 4936 10746
rect 4894 10704 4950 10713
rect 4894 10639 4950 10648
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4816 8634 4844 9318
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4816 6866 4844 7414
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4710 5808 4766 5817
rect 4710 5743 4766 5752
rect 4724 3414 4752 5743
rect 4894 5264 4950 5273
rect 4894 5199 4950 5208
rect 4908 4146 4936 5199
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4816 3534 4844 4082
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4724 3386 4844 3414
rect 4710 3088 4766 3097
rect 4710 3023 4712 3032
rect 4764 3023 4766 3032
rect 4712 2994 4764 3000
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4066 2615 4122 2624
rect 4252 2644 4304 2650
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 4080 1970 4108 2615
rect 4252 2586 4304 2592
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 4344 1964 4396 1970
rect 4344 1906 4396 1912
rect 4172 1601 4200 1906
rect 4158 1592 4214 1601
rect 4356 1562 4384 1906
rect 4712 1760 4764 1766
rect 4712 1702 4764 1708
rect 4158 1527 4214 1536
rect 4344 1556 4396 1562
rect 4344 1498 4396 1504
rect 3608 1352 3660 1358
rect 3606 1320 3608 1329
rect 4160 1352 4212 1358
rect 3660 1320 3662 1329
rect 3606 1255 3662 1264
rect 4066 1320 4122 1329
rect 4160 1294 4212 1300
rect 4066 1255 4068 1264
rect 4120 1255 4122 1264
rect 4068 1226 4120 1232
rect 570 1184 626 1193
rect 570 1119 626 1128
rect 3422 1184 3478 1193
rect 3422 1119 3478 1128
rect 3566 1116 3874 1125
rect 3566 1114 3572 1116
rect 3628 1114 3652 1116
rect 3708 1114 3732 1116
rect 3788 1114 3812 1116
rect 3868 1114 3874 1116
rect 3628 1062 3630 1114
rect 3810 1062 3812 1114
rect 3566 1060 3572 1062
rect 3628 1060 3652 1062
rect 3708 1060 3732 1062
rect 3788 1060 3812 1062
rect 3868 1060 3874 1062
rect 3566 1051 3874 1060
rect 386 912 442 921
rect 386 847 442 856
rect 4172 377 4200 1294
rect 4344 1216 4396 1222
rect 4344 1158 4396 1164
rect 4356 785 4384 1158
rect 4724 921 4752 1702
rect 4816 1358 4844 3386
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4908 3058 4936 3334
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4908 2582 4936 2994
rect 5000 2938 5028 7686
rect 5092 3738 5120 13262
rect 5276 12850 5304 14418
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5368 13920 5396 14282
rect 5460 14074 5488 14447
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5448 13932 5500 13938
rect 5368 13892 5448 13920
rect 5448 13874 5500 13880
rect 5460 13394 5488 13874
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5460 12434 5488 13330
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 12617 5580 13262
rect 5538 12608 5594 12617
rect 5538 12543 5594 12552
rect 5368 12406 5488 12434
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 8129 5212 11154
rect 5368 10674 5396 12406
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5170 8120 5226 8129
rect 5276 8090 5304 10406
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5368 8945 5396 9522
rect 5460 8974 5488 11018
rect 5448 8968 5500 8974
rect 5354 8936 5410 8945
rect 5448 8910 5500 8916
rect 5354 8871 5410 8880
rect 5170 8055 5226 8064
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5552 7857 5580 12038
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5644 10674 5672 10950
rect 5736 10742 5764 14962
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5920 13433 5948 13738
rect 5906 13424 5962 13433
rect 5906 13359 5962 13368
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5828 11830 5856 12718
rect 6012 12345 6040 16200
rect 6380 15706 6408 16759
rect 6458 16200 6514 17000
rect 16670 16960 16726 16969
rect 16670 16895 16726 16904
rect 13358 16824 13414 16833
rect 13358 16759 13414 16768
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6472 14482 6500 16200
rect 6826 16144 6882 16153
rect 6826 16079 6882 16088
rect 10874 16144 10930 16153
rect 10874 16079 10930 16088
rect 6840 15502 6868 16079
rect 7566 15804 7874 15813
rect 7566 15802 7572 15804
rect 7628 15802 7652 15804
rect 7708 15802 7732 15804
rect 7788 15802 7812 15804
rect 7868 15802 7874 15804
rect 7628 15750 7630 15802
rect 7810 15750 7812 15802
rect 7566 15748 7572 15750
rect 7628 15748 7652 15750
rect 7708 15748 7732 15750
rect 7788 15748 7812 15750
rect 7868 15748 7874 15750
rect 7566 15739 7874 15748
rect 6828 15496 6880 15502
rect 8392 15496 8444 15502
rect 6828 15438 6880 15444
rect 8114 15464 8170 15473
rect 7380 15428 7432 15434
rect 8392 15438 8444 15444
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 8114 15399 8116 15408
rect 7380 15370 7432 15376
rect 8168 15399 8170 15408
rect 8116 15370 8168 15376
rect 6644 15360 6696 15366
rect 6642 15328 6644 15337
rect 6696 15328 6698 15337
rect 6642 15263 6698 15272
rect 6550 15192 6606 15201
rect 6550 15127 6606 15136
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6564 12850 6592 15127
rect 7392 15094 7420 15370
rect 8404 15201 8432 15438
rect 8566 15260 8874 15269
rect 8566 15258 8572 15260
rect 8628 15258 8652 15260
rect 8708 15258 8732 15260
rect 8788 15258 8812 15260
rect 8868 15258 8874 15260
rect 8628 15206 8630 15258
rect 8810 15206 8812 15258
rect 8566 15204 8572 15206
rect 8628 15204 8652 15206
rect 8708 15204 8732 15206
rect 8788 15204 8812 15206
rect 8868 15204 8874 15206
rect 8390 15192 8446 15201
rect 8566 15195 8874 15204
rect 8390 15127 8446 15136
rect 7380 15088 7432 15094
rect 7300 15048 7380 15076
rect 7102 14376 7158 14385
rect 7102 14311 7158 14320
rect 7116 13938 7144 14311
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 5998 12336 6054 12345
rect 5998 12271 6054 12280
rect 6276 12232 6328 12238
rect 5906 12200 5962 12209
rect 6276 12174 6328 12180
rect 5906 12135 5908 12144
rect 5960 12135 5962 12144
rect 5908 12106 5960 12112
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5644 10169 5672 10610
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5722 10296 5778 10305
rect 5722 10231 5778 10240
rect 5630 10160 5686 10169
rect 5630 10095 5686 10104
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5644 8537 5672 8570
rect 5630 8528 5686 8537
rect 5630 8463 5686 8472
rect 5538 7848 5594 7857
rect 5264 7812 5316 7818
rect 5538 7783 5594 7792
rect 5264 7754 5316 7760
rect 5170 6896 5226 6905
rect 5170 6831 5226 6840
rect 5184 4826 5212 6831
rect 5276 5234 5304 7754
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5368 6254 5396 7482
rect 5538 7168 5594 7177
rect 5538 7103 5594 7112
rect 5552 6746 5580 7103
rect 5736 6882 5764 10231
rect 5828 10169 5856 10406
rect 5814 10160 5870 10169
rect 5814 10095 5870 10104
rect 5920 9994 5948 11494
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 6012 9761 6040 9998
rect 5998 9752 6054 9761
rect 5998 9687 6054 9696
rect 5814 9616 5870 9625
rect 5814 9551 5870 9560
rect 5828 9518 5856 9551
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5814 8800 5870 8809
rect 5814 8735 5870 8744
rect 5828 8498 5856 8735
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5906 8392 5962 8401
rect 5906 8327 5962 8336
rect 5736 6854 5856 6882
rect 5460 6718 5580 6746
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5722 6760 5778 6769
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5354 5944 5410 5953
rect 5354 5879 5410 5888
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5368 4978 5396 5879
rect 5276 4950 5396 4978
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5276 3670 5304 4950
rect 5354 4856 5410 4865
rect 5460 4826 5488 6718
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 5914 5580 6598
rect 5644 6458 5672 6734
rect 5722 6695 5778 6704
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5736 6186 5764 6695
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 5166 5580 5510
rect 5828 5234 5856 6854
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5354 4791 5410 4800
rect 5448 4820 5500 4826
rect 5368 4622 5396 4791
rect 5448 4762 5500 4768
rect 5828 4690 5856 5170
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5722 4584 5778 4593
rect 5722 4519 5778 4528
rect 5736 4146 5764 4519
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5460 3777 5488 3878
rect 5446 3768 5502 3777
rect 5446 3703 5502 3712
rect 5264 3664 5316 3670
rect 5644 3641 5672 4082
rect 5264 3606 5316 3612
rect 5630 3632 5686 3641
rect 5630 3567 5686 3576
rect 5078 3360 5134 3369
rect 5078 3295 5134 3304
rect 5092 3194 5120 3295
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5354 3088 5410 3097
rect 5354 3023 5356 3032
rect 5408 3023 5410 3032
rect 5356 2994 5408 3000
rect 5000 2910 5120 2938
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 4908 1970 4936 2518
rect 5000 2106 5028 2790
rect 4988 2100 5040 2106
rect 4988 2042 5040 2048
rect 4896 1964 4948 1970
rect 4896 1906 4948 1912
rect 5092 1358 5120 2910
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5460 2530 5488 2790
rect 5632 2576 5684 2582
rect 5630 2544 5632 2553
rect 5684 2544 5686 2553
rect 5460 2514 5580 2530
rect 5460 2508 5592 2514
rect 5460 2502 5540 2508
rect 5630 2479 5686 2488
rect 5540 2450 5592 2456
rect 5630 2408 5686 2417
rect 5630 2343 5686 2352
rect 5644 2106 5672 2343
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 5448 1964 5500 1970
rect 5448 1906 5500 1912
rect 5460 1601 5488 1906
rect 5446 1592 5502 1601
rect 5446 1527 5502 1536
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 5080 1352 5132 1358
rect 5080 1294 5132 1300
rect 5920 1222 5948 8327
rect 6104 6882 6132 10406
rect 6012 6854 6132 6882
rect 6012 6322 6040 6854
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6012 5642 6040 6258
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 6104 4826 6132 6734
rect 6196 5953 6224 10610
rect 6288 6905 6316 12174
rect 6564 11830 6592 12786
rect 6656 12442 6684 13194
rect 7300 13190 7328 15048
rect 7380 15030 7432 15036
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 7566 14716 7874 14725
rect 7566 14714 7572 14716
rect 7628 14714 7652 14716
rect 7708 14714 7732 14716
rect 7788 14714 7812 14716
rect 7868 14714 7874 14716
rect 7628 14662 7630 14714
rect 7810 14662 7812 14714
rect 7566 14660 7572 14662
rect 7628 14660 7652 14662
rect 7708 14660 7732 14662
rect 7788 14660 7812 14662
rect 7868 14660 7874 14662
rect 7566 14651 7874 14660
rect 8220 14414 8248 15030
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8956 14929 8984 14962
rect 8942 14920 8998 14929
rect 8942 14855 8998 14864
rect 8208 14408 8260 14414
rect 8260 14356 8340 14362
rect 8208 14350 8340 14356
rect 7380 14340 7432 14346
rect 8220 14334 8340 14350
rect 7380 14282 7432 14288
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12782 7328 13126
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6932 12306 6960 12718
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6918 12064 6974 12073
rect 6918 11999 6974 12008
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6380 8634 6408 9998
rect 6564 8838 6592 11766
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6656 9926 6684 11630
rect 6932 9994 6960 11999
rect 7300 11830 7328 12718
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 7300 11558 7328 11766
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7104 11144 7156 11150
rect 7010 11112 7066 11121
rect 7104 11086 7156 11092
rect 7194 11112 7250 11121
rect 7010 11047 7066 11056
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6828 9920 6880 9926
rect 7024 9897 7052 11047
rect 7010 9888 7066 9897
rect 6880 9868 6960 9874
rect 6828 9862 6960 9868
rect 6840 9846 6960 9862
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6380 7041 6408 7278
rect 6366 7032 6422 7041
rect 6366 6967 6422 6976
rect 6274 6896 6330 6905
rect 6472 6882 6500 8298
rect 6274 6831 6330 6840
rect 6380 6854 6500 6882
rect 6182 5944 6238 5953
rect 6182 5879 6238 5888
rect 6182 5672 6238 5681
rect 6182 5607 6238 5616
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6000 4752 6052 4758
rect 5998 4720 6000 4729
rect 6052 4720 6054 4729
rect 5998 4655 6054 4664
rect 6196 4622 6224 5607
rect 6184 4616 6236 4622
rect 5998 4584 6054 4593
rect 6184 4558 6236 4564
rect 5998 4519 6054 4528
rect 6012 3738 6040 4519
rect 6380 4146 6408 6854
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6472 5370 6500 6734
rect 6564 5817 6592 8774
rect 6932 8498 6960 9846
rect 7010 9823 7066 9832
rect 7024 9586 7052 9823
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7010 9344 7066 9353
rect 7010 9279 7066 9288
rect 7024 9042 7052 9279
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7024 8362 7052 8978
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 7116 8265 7144 11086
rect 7194 11047 7196 11056
rect 7248 11047 7250 11056
rect 7196 11018 7248 11024
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7102 8256 7158 8265
rect 7102 8191 7158 8200
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6828 6248 6880 6254
rect 6642 6216 6698 6225
rect 6828 6190 6880 6196
rect 6642 6151 6698 6160
rect 6550 5808 6606 5817
rect 6550 5743 6606 5752
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6564 5234 6592 5510
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6564 4214 6592 5170
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6656 4146 6684 6151
rect 6840 5352 6868 6190
rect 6932 5914 6960 7278
rect 7024 6322 7052 7686
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7116 7177 7144 7414
rect 7102 7168 7158 7177
rect 7102 7103 7158 7112
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6920 5364 6972 5370
rect 6840 5324 6920 5352
rect 6920 5306 6972 5312
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6748 4622 6776 5238
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6184 3936 6236 3942
rect 6182 3904 6184 3913
rect 6236 3904 6238 3913
rect 6182 3839 6238 3848
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 6380 3602 6408 4082
rect 6840 3618 6868 4966
rect 7116 4282 7144 6666
rect 7208 6089 7236 10678
rect 7392 9654 7420 14282
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 8022 13968 8078 13977
rect 7566 13628 7874 13637
rect 7566 13626 7572 13628
rect 7628 13626 7652 13628
rect 7708 13626 7732 13628
rect 7788 13626 7812 13628
rect 7868 13626 7874 13628
rect 7628 13574 7630 13626
rect 7810 13574 7812 13626
rect 7566 13572 7572 13574
rect 7628 13572 7652 13574
rect 7708 13572 7732 13574
rect 7788 13572 7812 13574
rect 7868 13572 7874 13574
rect 7566 13563 7874 13572
rect 7566 12540 7874 12549
rect 7566 12538 7572 12540
rect 7628 12538 7652 12540
rect 7708 12538 7732 12540
rect 7788 12538 7812 12540
rect 7868 12538 7874 12540
rect 7628 12486 7630 12538
rect 7810 12486 7812 12538
rect 7566 12484 7572 12486
rect 7628 12484 7652 12486
rect 7708 12484 7732 12486
rect 7788 12484 7812 12486
rect 7868 12484 7874 12486
rect 7566 12475 7874 12484
rect 7566 11452 7874 11461
rect 7566 11450 7572 11452
rect 7628 11450 7652 11452
rect 7708 11450 7732 11452
rect 7788 11450 7812 11452
rect 7868 11450 7874 11452
rect 7628 11398 7630 11450
rect 7810 11398 7812 11450
rect 7566 11396 7572 11398
rect 7628 11396 7652 11398
rect 7708 11396 7732 11398
rect 7788 11396 7812 11398
rect 7868 11396 7874 11398
rect 7566 11387 7874 11396
rect 7944 10606 7972 13942
rect 8022 13903 8078 13912
rect 8036 10810 8064 13903
rect 8208 13184 8260 13190
rect 8114 13152 8170 13161
rect 8208 13126 8260 13132
rect 8114 13087 8170 13096
rect 8128 12434 8156 13087
rect 8220 12889 8248 13126
rect 8312 12986 8340 14334
rect 8392 14340 8444 14346
rect 8392 14282 8444 14288
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8206 12880 8262 12889
rect 8206 12815 8262 12824
rect 8128 12406 8248 12434
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8128 11898 8156 12242
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8220 10962 8248 12406
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8128 10934 8248 10962
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7566 10364 7874 10373
rect 7566 10362 7572 10364
rect 7628 10362 7652 10364
rect 7708 10362 7732 10364
rect 7788 10362 7812 10364
rect 7868 10362 7874 10364
rect 7628 10310 7630 10362
rect 7810 10310 7812 10362
rect 7566 10308 7572 10310
rect 7628 10308 7652 10310
rect 7708 10308 7732 10310
rect 7788 10308 7812 10310
rect 7868 10308 7874 10310
rect 7566 10299 7874 10308
rect 8022 10024 8078 10033
rect 8022 9959 8078 9968
rect 8036 9926 8064 9959
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7194 6080 7250 6089
rect 7194 6015 7250 6024
rect 7194 5128 7250 5137
rect 7194 5063 7250 5072
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7010 3632 7066 3641
rect 6368 3596 6420 3602
rect 6840 3590 6960 3618
rect 6368 3538 6420 3544
rect 5998 3496 6054 3505
rect 5998 3431 6054 3440
rect 6012 3058 6040 3431
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 6380 2774 6408 3538
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6288 2746 6408 2774
rect 6090 2544 6146 2553
rect 6090 2479 6146 2488
rect 6104 1970 6132 2479
rect 6288 2446 6316 2746
rect 6276 2440 6328 2446
rect 6644 2440 6696 2446
rect 6276 2382 6328 2388
rect 6564 2388 6644 2394
rect 6564 2382 6696 2388
rect 6288 2258 6316 2382
rect 6196 2230 6316 2258
rect 6564 2366 6684 2382
rect 6196 1970 6224 2230
rect 6276 2100 6328 2106
rect 6276 2042 6328 2048
rect 6288 2009 6316 2042
rect 6274 2000 6330 2009
rect 6092 1964 6144 1970
rect 6092 1906 6144 1912
rect 6184 1964 6236 1970
rect 6274 1935 6330 1944
rect 6184 1906 6236 1912
rect 6196 1358 6224 1906
rect 6564 1737 6592 2366
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6550 1728 6606 1737
rect 6550 1663 6606 1672
rect 6184 1352 6236 1358
rect 6184 1294 6236 1300
rect 4896 1216 4948 1222
rect 4896 1158 4948 1164
rect 5908 1216 5960 1222
rect 5908 1158 5960 1164
rect 4908 921 4936 1158
rect 4710 912 4766 921
rect 4710 847 4766 856
rect 4894 912 4950 921
rect 4894 847 4950 856
rect 4342 776 4398 785
rect 4342 711 4398 720
rect 6656 513 6684 2246
rect 6748 1970 6776 2246
rect 6840 1986 6868 3470
rect 6932 3126 6960 3590
rect 7010 3567 7066 3576
rect 7024 3534 7052 3567
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7208 3210 7236 5063
rect 7300 4865 7328 8910
rect 7392 7886 7420 9590
rect 7566 9276 7874 9285
rect 7566 9274 7572 9276
rect 7628 9274 7652 9276
rect 7708 9274 7732 9276
rect 7788 9274 7812 9276
rect 7868 9274 7874 9276
rect 7628 9222 7630 9274
rect 7810 9222 7812 9274
rect 7566 9220 7572 9222
rect 7628 9220 7652 9222
rect 7708 9220 7732 9222
rect 7788 9220 7812 9222
rect 7868 9220 7874 9222
rect 7566 9211 7874 9220
rect 8022 9208 8078 9217
rect 8022 9143 8078 9152
rect 8036 8809 8064 9143
rect 8022 8800 8078 8809
rect 8022 8735 8078 8744
rect 7566 8188 7874 8197
rect 7566 8186 7572 8188
rect 7628 8186 7652 8188
rect 7708 8186 7732 8188
rect 7788 8186 7812 8188
rect 7868 8186 7874 8188
rect 7628 8134 7630 8186
rect 7810 8134 7812 8186
rect 7566 8132 7572 8134
rect 7628 8132 7652 8134
rect 7708 8132 7732 8134
rect 7788 8132 7812 8134
rect 7868 8132 7874 8134
rect 7566 8123 7874 8132
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8036 7546 8064 7822
rect 8128 7818 8156 10934
rect 8312 10674 8340 12038
rect 8404 10674 8432 14282
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8496 13938 8524 14214
rect 8566 14172 8874 14181
rect 8566 14170 8572 14172
rect 8628 14170 8652 14172
rect 8708 14170 8732 14172
rect 8788 14170 8812 14172
rect 8868 14170 8874 14172
rect 8628 14118 8630 14170
rect 8810 14118 8812 14170
rect 8566 14116 8572 14118
rect 8628 14116 8652 14118
rect 8708 14116 8732 14118
rect 8788 14116 8812 14118
rect 8868 14116 8874 14118
rect 8566 14107 8874 14116
rect 8942 13968 8998 13977
rect 8484 13932 8536 13938
rect 8942 13903 8944 13912
rect 8484 13874 8536 13880
rect 8996 13903 8998 13912
rect 8944 13874 8996 13880
rect 8566 13084 8874 13093
rect 8566 13082 8572 13084
rect 8628 13082 8652 13084
rect 8708 13082 8732 13084
rect 8788 13082 8812 13084
rect 8868 13082 8874 13084
rect 8628 13030 8630 13082
rect 8810 13030 8812 13082
rect 8566 13028 8572 13030
rect 8628 13028 8652 13030
rect 8708 13028 8732 13030
rect 8788 13028 8812 13030
rect 8868 13028 8874 13030
rect 8566 13019 8874 13028
rect 8942 12336 8998 12345
rect 8942 12271 8998 12280
rect 8956 12238 8984 12271
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8496 11082 8524 12106
rect 8566 11996 8874 12005
rect 8566 11994 8572 11996
rect 8628 11994 8652 11996
rect 8708 11994 8732 11996
rect 8788 11994 8812 11996
rect 8868 11994 8874 11996
rect 8628 11942 8630 11994
rect 8810 11942 8812 11994
rect 8566 11940 8572 11942
rect 8628 11940 8652 11942
rect 8708 11940 8732 11942
rect 8788 11940 8812 11942
rect 8868 11940 8874 11942
rect 8566 11931 8874 11940
rect 9048 11898 9076 15438
rect 9128 15360 9180 15366
rect 9126 15328 9128 15337
rect 9180 15328 9182 15337
rect 9126 15263 9182 15272
rect 10690 14920 10746 14929
rect 10690 14855 10746 14864
rect 10704 14482 10732 14855
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 10322 14376 10378 14385
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9324 14113 9352 14214
rect 9310 14104 9366 14113
rect 9310 14039 9366 14048
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8852 11824 8904 11830
rect 8850 11792 8852 11801
rect 8904 11792 8906 11801
rect 8760 11756 8812 11762
rect 8850 11727 8906 11736
rect 8944 11756 8996 11762
rect 8760 11698 8812 11704
rect 8944 11698 8996 11704
rect 8772 11393 8800 11698
rect 8758 11384 8814 11393
rect 8758 11319 8814 11328
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8566 10908 8874 10917
rect 8566 10906 8572 10908
rect 8628 10906 8652 10908
rect 8708 10906 8732 10908
rect 8788 10906 8812 10908
rect 8868 10906 8874 10908
rect 8628 10854 8630 10906
rect 8810 10854 8812 10906
rect 8566 10852 8572 10854
rect 8628 10852 8652 10854
rect 8708 10852 8732 10854
rect 8788 10852 8812 10854
rect 8868 10852 8874 10854
rect 8566 10843 8874 10852
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8220 9897 8248 9930
rect 8206 9888 8262 9897
rect 8206 9823 8262 9832
rect 8298 9752 8354 9761
rect 8298 9687 8354 9696
rect 8208 8424 8260 8430
rect 8206 8392 8208 8401
rect 8260 8392 8262 8401
rect 8206 8327 8262 8336
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7566 7100 7874 7109
rect 7566 7098 7572 7100
rect 7628 7098 7652 7100
rect 7708 7098 7732 7100
rect 7788 7098 7812 7100
rect 7868 7098 7874 7100
rect 7628 7046 7630 7098
rect 7810 7046 7812 7098
rect 7566 7044 7572 7046
rect 7628 7044 7652 7046
rect 7708 7044 7732 7046
rect 7788 7044 7812 7046
rect 7868 7044 7874 7046
rect 7566 7035 7874 7044
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7286 4856 7342 4865
rect 7392 4826 7420 6326
rect 7286 4791 7342 4800
rect 7380 4820 7432 4826
rect 7300 4706 7328 4791
rect 7380 4762 7432 4768
rect 7300 4678 7420 4706
rect 7392 4622 7420 4678
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7392 4282 7420 4558
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7116 3194 7236 3210
rect 7104 3188 7236 3194
rect 7156 3182 7236 3188
rect 7104 3130 7156 3136
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 7300 3058 7328 3878
rect 7484 3194 7512 6734
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7566 6012 7874 6021
rect 7566 6010 7572 6012
rect 7628 6010 7652 6012
rect 7708 6010 7732 6012
rect 7788 6010 7812 6012
rect 7868 6010 7874 6012
rect 7628 5958 7630 6010
rect 7810 5958 7812 6010
rect 7566 5956 7572 5958
rect 7628 5956 7652 5958
rect 7708 5956 7732 5958
rect 7788 5956 7812 5958
rect 7868 5956 7874 5958
rect 7566 5947 7874 5956
rect 7944 5574 7972 6598
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7566 4924 7874 4933
rect 7566 4922 7572 4924
rect 7628 4922 7652 4924
rect 7708 4922 7732 4924
rect 7788 4922 7812 4924
rect 7868 4922 7874 4924
rect 7628 4870 7630 4922
rect 7810 4870 7812 4922
rect 7566 4868 7572 4870
rect 7628 4868 7652 4870
rect 7708 4868 7732 4870
rect 7788 4868 7812 4870
rect 7868 4868 7874 4870
rect 7566 4859 7874 4868
rect 7566 3836 7874 3845
rect 7566 3834 7572 3836
rect 7628 3834 7652 3836
rect 7708 3834 7732 3836
rect 7788 3834 7812 3836
rect 7868 3834 7874 3836
rect 7628 3782 7630 3834
rect 7810 3782 7812 3834
rect 7566 3780 7572 3782
rect 7628 3780 7652 3782
rect 7708 3780 7732 3782
rect 7788 3780 7812 3782
rect 7868 3780 7874 3782
rect 7566 3771 7874 3780
rect 7944 3482 7972 5170
rect 7852 3454 7972 3482
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7852 2938 7880 3454
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 3074 7972 3334
rect 8036 3194 8064 7346
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8128 4690 8156 6734
rect 8206 6080 8262 6089
rect 8206 6015 8262 6024
rect 8220 5710 8248 6015
rect 8312 5914 8340 9687
rect 8404 6905 8432 10610
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8390 6896 8446 6905
rect 8390 6831 8446 6840
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8208 4480 8260 4486
rect 8206 4448 8208 4457
rect 8260 4448 8262 4457
rect 8206 4383 8262 4392
rect 8312 4162 8340 5714
rect 8404 5710 8432 6831
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8220 4134 8340 4162
rect 8220 3942 8248 4134
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8206 3768 8262 3777
rect 8206 3703 8262 3712
rect 8220 3534 8248 3703
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8404 3482 8432 5510
rect 8496 4826 8524 9998
rect 8680 9926 8708 10746
rect 8956 10266 8984 11698
rect 9140 11370 9168 13262
rect 9310 12608 9366 12617
rect 9310 12543 9366 12552
rect 9140 11342 9260 11370
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8566 9820 8874 9829
rect 8566 9818 8572 9820
rect 8628 9818 8652 9820
rect 8708 9818 8732 9820
rect 8788 9818 8812 9820
rect 8868 9818 8874 9820
rect 8628 9766 8630 9818
rect 8810 9766 8812 9818
rect 8566 9764 8572 9766
rect 8628 9764 8652 9766
rect 8708 9764 8732 9766
rect 8788 9764 8812 9766
rect 8868 9764 8874 9766
rect 8566 9755 8874 9764
rect 8942 9616 8998 9625
rect 9048 9602 9076 11086
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9140 10266 9168 10746
rect 9232 10713 9260 11342
rect 9218 10704 9274 10713
rect 9218 10639 9274 10648
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9128 9920 9180 9926
rect 9126 9888 9128 9897
rect 9180 9888 9182 9897
rect 9126 9823 9182 9832
rect 8998 9574 9076 9602
rect 8942 9551 8998 9560
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 8974 9076 9318
rect 9036 8968 9088 8974
rect 8942 8936 8998 8945
rect 9036 8910 9088 8916
rect 8942 8871 8998 8880
rect 8566 8732 8874 8741
rect 8566 8730 8572 8732
rect 8628 8730 8652 8732
rect 8708 8730 8732 8732
rect 8788 8730 8812 8732
rect 8868 8730 8874 8732
rect 8628 8678 8630 8730
rect 8810 8678 8812 8730
rect 8566 8676 8572 8678
rect 8628 8676 8652 8678
rect 8708 8676 8732 8678
rect 8788 8676 8812 8678
rect 8868 8676 8874 8678
rect 8566 8667 8874 8676
rect 8566 7644 8874 7653
rect 8566 7642 8572 7644
rect 8628 7642 8652 7644
rect 8708 7642 8732 7644
rect 8788 7642 8812 7644
rect 8868 7642 8874 7644
rect 8628 7590 8630 7642
rect 8810 7590 8812 7642
rect 8566 7588 8572 7590
rect 8628 7588 8652 7590
rect 8708 7588 8732 7590
rect 8788 7588 8812 7590
rect 8868 7588 8874 7590
rect 8566 7579 8874 7588
rect 8956 7546 8984 8871
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9140 8566 9168 8774
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 9048 7426 9076 7822
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 8864 7398 9076 7426
rect 8864 6730 8892 7398
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8566 6556 8874 6565
rect 8566 6554 8572 6556
rect 8628 6554 8652 6556
rect 8708 6554 8732 6556
rect 8788 6554 8812 6556
rect 8868 6554 8874 6556
rect 8628 6502 8630 6554
rect 8810 6502 8812 6554
rect 8566 6500 8572 6502
rect 8628 6500 8652 6502
rect 8708 6500 8732 6502
rect 8788 6500 8812 6502
rect 8868 6500 8874 6502
rect 8566 6491 8874 6500
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8864 5681 8892 6054
rect 8850 5672 8906 5681
rect 8850 5607 8906 5616
rect 8566 5468 8874 5477
rect 8566 5466 8572 5468
rect 8628 5466 8652 5468
rect 8708 5466 8732 5468
rect 8788 5466 8812 5468
rect 8868 5466 8874 5468
rect 8628 5414 8630 5466
rect 8810 5414 8812 5466
rect 8566 5412 8572 5414
rect 8628 5412 8652 5414
rect 8708 5412 8732 5414
rect 8788 5412 8812 5414
rect 8868 5412 8874 5414
rect 8566 5403 8874 5412
rect 8574 4992 8630 5001
rect 8574 4927 8630 4936
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8588 4622 8616 4927
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8566 4380 8874 4389
rect 8566 4378 8572 4380
rect 8628 4378 8652 4380
rect 8708 4378 8732 4380
rect 8788 4378 8812 4380
rect 8868 4378 8874 4380
rect 8628 4326 8630 4378
rect 8810 4326 8812 4378
rect 8566 4324 8572 4326
rect 8628 4324 8652 4326
rect 8708 4324 8732 4326
rect 8788 4324 8812 4326
rect 8868 4324 8874 4326
rect 8566 4315 8874 4324
rect 8956 3534 8984 7142
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 5658 9076 6598
rect 9140 6225 9168 7686
rect 9126 6216 9182 6225
rect 9126 6151 9182 6160
rect 9232 5794 9260 7686
rect 9324 6798 9352 12543
rect 9416 12170 9444 14282
rect 9508 12594 9536 14350
rect 10322 14311 10324 14320
rect 10376 14311 10378 14320
rect 10324 14282 10376 14288
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9508 12566 9674 12594
rect 9646 12434 9674 12566
rect 9784 12434 9812 14010
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 9646 12406 9720 12434
rect 9784 12406 10088 12434
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9692 10849 9720 12406
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9678 10840 9734 10849
rect 9678 10775 9734 10784
rect 9494 10568 9550 10577
rect 9494 10503 9550 10512
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9140 5778 9260 5794
rect 9128 5772 9260 5778
rect 9180 5766 9260 5772
rect 9128 5714 9180 5720
rect 9220 5704 9272 5710
rect 9048 5630 9168 5658
rect 9220 5646 9272 5652
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 8944 3528 8996 3534
rect 8404 3454 8524 3482
rect 8944 3470 8996 3476
rect 8116 3392 8168 3398
rect 8392 3392 8444 3398
rect 8116 3334 8168 3340
rect 8390 3360 8392 3369
rect 8444 3360 8446 3369
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7944 3046 8064 3074
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7208 2666 7236 2858
rect 7116 2638 7236 2666
rect 7116 2378 7144 2638
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 6840 1970 7052 1986
rect 6736 1964 6788 1970
rect 6840 1964 7064 1970
rect 6840 1958 7012 1964
rect 6736 1906 6788 1912
rect 7012 1906 7064 1912
rect 6828 1760 6880 1766
rect 6828 1702 6880 1708
rect 6840 1465 6868 1702
rect 6826 1456 6882 1465
rect 7484 1442 7512 2926
rect 7852 2910 7972 2938
rect 7566 2748 7874 2757
rect 7566 2746 7572 2748
rect 7628 2746 7652 2748
rect 7708 2746 7732 2748
rect 7788 2746 7812 2748
rect 7868 2746 7874 2748
rect 7628 2694 7630 2746
rect 7810 2694 7812 2746
rect 7566 2692 7572 2694
rect 7628 2692 7652 2694
rect 7708 2692 7732 2694
rect 7788 2692 7812 2694
rect 7868 2692 7874 2694
rect 7566 2683 7874 2692
rect 7944 2514 7972 2910
rect 8036 2825 8064 3046
rect 8022 2816 8078 2825
rect 8022 2751 8078 2760
rect 8022 2680 8078 2689
rect 8022 2615 8078 2624
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8036 2106 8064 2615
rect 8024 2100 8076 2106
rect 8024 2042 8076 2048
rect 8128 2038 8156 3334
rect 8390 3295 8446 3304
rect 8496 3058 8524 3454
rect 8566 3292 8874 3301
rect 8566 3290 8572 3292
rect 8628 3290 8652 3292
rect 8708 3290 8732 3292
rect 8788 3290 8812 3292
rect 8868 3290 8874 3292
rect 8628 3238 8630 3290
rect 8810 3238 8812 3290
rect 8566 3236 8572 3238
rect 8628 3236 8652 3238
rect 8708 3236 8732 3238
rect 8788 3236 8812 3238
rect 8868 3236 8874 3238
rect 8566 3227 8874 3236
rect 9048 3058 9076 5510
rect 9140 4146 9168 5630
rect 9232 5302 9260 5646
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9218 5128 9274 5137
rect 9218 5063 9274 5072
rect 9232 4826 9260 5063
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9220 3936 9272 3942
rect 9218 3904 9220 3913
rect 9272 3904 9274 3913
rect 9218 3839 9274 3848
rect 9218 3224 9274 3233
rect 9218 3159 9220 3168
rect 9272 3159 9274 3168
rect 9220 3130 9272 3136
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8208 2440 8260 2446
rect 8312 2428 8340 2790
rect 9232 2650 9260 2994
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 8482 2544 8538 2553
rect 8482 2479 8538 2488
rect 8260 2400 8340 2428
rect 8208 2382 8260 2388
rect 8496 2106 8524 2479
rect 9324 2446 9352 6598
rect 9416 4622 9444 10066
rect 9508 8634 9536 10503
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9600 8498 9628 8774
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9508 7410 9536 8026
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9508 3126 9536 5578
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 8566 2204 8874 2213
rect 8566 2202 8572 2204
rect 8628 2202 8652 2204
rect 8708 2202 8732 2204
rect 8788 2202 8812 2204
rect 8868 2202 8874 2204
rect 8628 2150 8630 2202
rect 8810 2150 8812 2202
rect 8566 2148 8572 2150
rect 8628 2148 8652 2150
rect 8708 2148 8732 2150
rect 8788 2148 8812 2150
rect 8868 2148 8874 2150
rect 8566 2139 8874 2148
rect 8484 2100 8536 2106
rect 8484 2042 8536 2048
rect 8116 2032 8168 2038
rect 8116 1974 8168 1980
rect 9600 1970 9628 8434
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9678 5808 9734 5817
rect 9678 5743 9734 5752
rect 9692 4593 9720 5743
rect 9678 4584 9734 4593
rect 9678 4519 9734 4528
rect 9784 2582 9812 6258
rect 9862 5536 9918 5545
rect 9862 5471 9918 5480
rect 9876 3398 9904 5471
rect 9968 4486 9996 12038
rect 10060 9217 10088 12406
rect 10152 10266 10180 12582
rect 10888 12374 10916 16079
rect 11886 16008 11942 16017
rect 11886 15943 11942 15952
rect 11058 15600 11114 15609
rect 11058 15535 11114 15544
rect 11072 14657 11100 15535
rect 11702 15328 11758 15337
rect 11702 15263 11758 15272
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11058 14648 11114 14657
rect 11058 14583 11114 14592
rect 11058 14104 11114 14113
rect 11058 14039 11114 14048
rect 11072 12617 11100 14039
rect 11058 12608 11114 12617
rect 11058 12543 11114 12552
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 11440 11830 11468 14758
rect 11610 12744 11666 12753
rect 11610 12679 11666 12688
rect 11624 11898 11652 12679
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11716 11150 11744 15263
rect 11794 12880 11850 12889
rect 11794 12815 11850 12824
rect 11808 11937 11836 12815
rect 11794 11928 11850 11937
rect 11794 11863 11850 11872
rect 11900 11801 11928 15943
rect 12898 14512 12954 14521
rect 12898 14447 12954 14456
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 12176 12918 12204 13194
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 12714 12064 12770 12073
rect 12714 11999 12770 12008
rect 11886 11792 11942 11801
rect 11886 11727 11942 11736
rect 12530 11384 12586 11393
rect 12530 11319 12586 11328
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 12438 10432 12494 10441
rect 12438 10367 12494 10376
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 11704 9784 11756 9790
rect 11704 9726 11756 9732
rect 11716 9489 11744 9726
rect 11702 9480 11758 9489
rect 11702 9415 11758 9424
rect 10046 9208 10102 9217
rect 10046 9143 10102 9152
rect 10060 5234 10088 9143
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10520 6089 10548 8366
rect 11794 8256 11850 8265
rect 11794 8191 11850 8200
rect 10784 7132 10836 7138
rect 10784 7074 10836 7080
rect 10506 6080 10562 6089
rect 10506 6015 10562 6024
rect 10322 5400 10378 5409
rect 10322 5335 10378 5344
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 8484 1896 8536 1902
rect 8482 1864 8484 1873
rect 8668 1896 8720 1902
rect 8536 1864 8538 1873
rect 8668 1838 8720 1844
rect 8482 1799 8538 1808
rect 8680 1737 8708 1838
rect 10336 1737 10364 5335
rect 10690 3496 10746 3505
rect 10690 3431 10746 3440
rect 10704 2417 10732 3431
rect 10690 2408 10746 2417
rect 10690 2343 10746 2352
rect 8666 1728 8722 1737
rect 7566 1660 7874 1669
rect 8666 1663 8722 1672
rect 10322 1728 10378 1737
rect 10322 1663 10378 1672
rect 7566 1658 7572 1660
rect 7628 1658 7652 1660
rect 7708 1658 7732 1660
rect 7788 1658 7812 1660
rect 7868 1658 7874 1660
rect 7628 1606 7630 1658
rect 7810 1606 7812 1658
rect 7566 1604 7572 1606
rect 7628 1604 7652 1606
rect 7708 1604 7732 1606
rect 7788 1604 7812 1606
rect 7868 1604 7874 1606
rect 7566 1595 7874 1604
rect 6826 1391 6882 1400
rect 7116 1414 7512 1442
rect 6736 1352 6788 1358
rect 7116 1306 7144 1414
rect 7380 1352 7432 1358
rect 6736 1294 6788 1300
rect 6748 649 6776 1294
rect 6840 1290 7144 1306
rect 6828 1284 7144 1290
rect 6880 1278 7144 1284
rect 7378 1320 7380 1329
rect 10796 1329 10824 7074
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10888 3097 10916 6938
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11058 5672 11114 5681
rect 11058 5607 11114 5616
rect 11072 5273 11100 5607
rect 11058 5264 11114 5273
rect 11058 5199 11114 5208
rect 11058 4448 11114 4457
rect 11058 4383 11114 4392
rect 11072 3641 11100 4383
rect 11058 3632 11114 3641
rect 11058 3567 11114 3576
rect 10874 3088 10930 3097
rect 10874 3023 10930 3032
rect 7432 1320 7434 1329
rect 7378 1255 7434 1264
rect 10782 1320 10838 1329
rect 10782 1255 10838 1264
rect 6828 1226 6880 1232
rect 7288 1216 7340 1222
rect 7288 1158 7340 1164
rect 7300 785 7328 1158
rect 8566 1116 8874 1125
rect 8566 1114 8572 1116
rect 8628 1114 8652 1116
rect 8708 1114 8732 1116
rect 8788 1114 8812 1116
rect 8868 1114 8874 1116
rect 8628 1062 8630 1114
rect 8810 1062 8812 1114
rect 8566 1060 8572 1062
rect 8628 1060 8652 1062
rect 8708 1060 8732 1062
rect 8788 1060 8812 1062
rect 8868 1060 8874 1062
rect 8566 1051 8874 1060
rect 7102 776 7158 785
rect 7102 711 7158 720
rect 7286 776 7342 785
rect 7286 711 7342 720
rect 6734 640 6790 649
rect 6734 575 6790 584
rect 7116 513 7144 711
rect 6642 504 6698 513
rect 6642 439 6698 448
rect 6918 504 6974 513
rect 6918 439 6974 448
rect 7102 504 7158 513
rect 7102 439 7158 448
rect 4158 368 4214 377
rect 4158 303 4214 312
rect 6932 241 6960 439
rect 11164 241 11192 6802
rect 11808 6769 11836 8191
rect 11886 7032 11942 7041
rect 11886 6967 11942 6976
rect 11794 6760 11850 6769
rect 11794 6695 11850 6704
rect 11242 6624 11298 6633
rect 11242 6559 11298 6568
rect 11256 3738 11284 6559
rect 11334 5264 11390 5273
rect 11334 5199 11390 5208
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11242 3632 11298 3641
rect 11242 3567 11298 3576
rect 11256 2922 11284 3567
rect 11348 2990 11376 5199
rect 11900 4729 11928 6967
rect 12346 6216 12402 6225
rect 12346 6151 12402 6160
rect 11886 4720 11942 4729
rect 11886 4655 11942 4664
rect 11794 4584 11850 4593
rect 11794 4519 11850 4528
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11808 1873 11836 4519
rect 11794 1864 11850 1873
rect 11794 1799 11850 1808
rect 12360 1465 12388 6151
rect 12452 5001 12480 10367
rect 12544 5273 12572 11319
rect 12622 10024 12678 10033
rect 12622 9959 12678 9968
rect 12530 5264 12586 5273
rect 12530 5199 12586 5208
rect 12438 4992 12494 5001
rect 12438 4927 12494 4936
rect 12636 3777 12664 9959
rect 12728 5545 12756 11999
rect 12806 11656 12862 11665
rect 12806 11591 12862 11600
rect 12714 5536 12770 5545
rect 12714 5471 12770 5480
rect 12622 3768 12678 3777
rect 12622 3703 12678 3712
rect 12820 3641 12848 11591
rect 12912 6225 12940 14447
rect 13174 12608 13230 12617
rect 13174 12543 13176 12552
rect 13228 12543 13230 12552
rect 13176 12514 13228 12520
rect 13372 12481 13400 16759
rect 15842 16688 15898 16697
rect 15842 16623 15898 16632
rect 13726 15464 13782 15473
rect 13726 15399 13782 15408
rect 13740 13977 13768 15399
rect 13818 14784 13874 14793
rect 13818 14719 13820 14728
rect 13872 14719 13874 14728
rect 13820 14690 13872 14696
rect 14096 14340 14148 14346
rect 14096 14282 14148 14288
rect 13542 13968 13598 13977
rect 13542 13903 13598 13912
rect 13726 13968 13782 13977
rect 13726 13903 13782 13912
rect 13450 13832 13506 13841
rect 13450 13767 13506 13776
rect 13358 12472 13414 12481
rect 13358 12407 13414 12416
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13372 11121 13400 11154
rect 13358 11112 13414 11121
rect 13358 11047 13414 11056
rect 13082 9888 13138 9897
rect 13082 9823 13138 9832
rect 12990 8392 13046 8401
rect 12990 8327 13046 8336
rect 12898 6216 12954 6225
rect 12898 6151 12954 6160
rect 13004 5001 13032 8327
rect 13096 6254 13124 9823
rect 13266 7440 13322 7449
rect 13266 7375 13322 7384
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 12990 4992 13046 5001
rect 12990 4927 13046 4936
rect 12806 3632 12862 3641
rect 12806 3567 12862 3576
rect 13188 2961 13216 6666
rect 13280 3913 13308 7375
rect 13358 6216 13414 6225
rect 13358 6151 13414 6160
rect 13266 3904 13322 3913
rect 13266 3839 13322 3848
rect 13174 2952 13230 2961
rect 13174 2887 13230 2896
rect 13372 2514 13400 6151
rect 13464 5817 13492 13767
rect 13450 5808 13506 5817
rect 13450 5743 13506 5752
rect 13556 5681 13584 13903
rect 13634 13424 13690 13433
rect 13634 13359 13690 13368
rect 13648 6730 13676 13359
rect 13818 13152 13874 13161
rect 13818 13087 13820 13096
rect 13872 13087 13874 13096
rect 13820 13058 13872 13064
rect 13912 12572 13964 12578
rect 13912 12514 13964 12520
rect 13924 12434 13952 12514
rect 13924 12406 14044 12434
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13740 10713 13768 11766
rect 13820 11144 13872 11150
rect 13818 11112 13820 11121
rect 13872 11112 13874 11121
rect 13818 11047 13874 11056
rect 13818 10840 13874 10849
rect 13874 10798 13952 10826
rect 13818 10775 13874 10784
rect 13726 10704 13782 10713
rect 13726 10639 13782 10648
rect 13820 9920 13872 9926
rect 13818 9888 13820 9897
rect 13872 9888 13874 9897
rect 13818 9823 13874 9832
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13832 9489 13860 9658
rect 13818 9480 13874 9489
rect 13818 9415 13874 9424
rect 13820 9240 13872 9246
rect 13820 9182 13872 9188
rect 13832 9081 13860 9182
rect 13818 9072 13874 9081
rect 13818 9007 13874 9016
rect 13726 7848 13782 7857
rect 13726 7783 13782 7792
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13542 5672 13598 5681
rect 13542 5607 13598 5616
rect 13740 5137 13768 7783
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13832 6361 13860 6394
rect 13818 6352 13874 6361
rect 13818 6287 13874 6296
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13832 5817 13860 6122
rect 13818 5808 13874 5817
rect 13818 5743 13874 5752
rect 13832 5642 13860 5743
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13726 5128 13782 5137
rect 13726 5063 13782 5072
rect 13820 4888 13872 4894
rect 13818 4856 13820 4865
rect 13872 4856 13874 4865
rect 13818 4791 13874 4800
rect 13924 4570 13952 10798
rect 13740 4542 13952 4570
rect 13740 4457 13768 4542
rect 13726 4448 13782 4457
rect 13726 4383 13782 4392
rect 14016 3369 14044 12406
rect 14108 4894 14136 14282
rect 15152 13560 15208 13569
rect 15208 13518 15332 13546
rect 15152 13495 15208 13504
rect 15304 12442 15332 13518
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15028 8242 15056 12378
rect 15152 12336 15208 12345
rect 15488 12322 15516 12786
rect 15208 12294 15516 12322
rect 15152 12271 15208 12280
rect 15488 11626 15516 12294
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15152 11520 15208 11529
rect 15208 11478 15516 11506
rect 15152 11455 15208 11464
rect 15292 11416 15344 11422
rect 15292 11358 15344 11364
rect 15304 10418 15332 11358
rect 15488 11150 15516 11478
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15384 10940 15436 10946
rect 15384 10882 15436 10888
rect 15166 10390 15332 10418
rect 15166 10305 15194 10390
rect 15152 10296 15208 10305
rect 15152 10231 15208 10240
rect 15108 9920 15160 9926
rect 15160 9868 15240 9874
rect 15108 9862 15240 9868
rect 15120 9846 15240 9862
rect 15108 9716 15160 9722
rect 15212 9704 15240 9846
rect 15212 9676 15332 9704
rect 15108 9658 15160 9664
rect 15120 9568 15148 9658
rect 15200 9580 15252 9586
rect 15120 9540 15200 9568
rect 15200 9522 15252 9528
rect 15304 8838 15332 9676
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15028 8214 15332 8242
rect 14096 4888 14148 4894
rect 14096 4830 14148 4836
rect 14554 4312 14610 4321
rect 14554 4247 14610 4256
rect 14002 3360 14058 3369
rect 14002 3295 14058 3304
rect 14568 2825 14596 4247
rect 14554 2816 14610 2825
rect 14554 2751 14610 2760
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 15304 2009 15332 8214
rect 15396 7138 15424 10882
rect 15488 9586 15516 10950
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15580 9246 15608 13126
rect 15660 13116 15712 13122
rect 15660 13058 15712 13064
rect 15672 11286 15700 13058
rect 15752 11620 15804 11626
rect 15752 11562 15804 11568
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15568 9240 15620 9246
rect 15568 9182 15620 9188
rect 15384 7132 15436 7138
rect 15384 7074 15436 7080
rect 15672 6458 15700 11086
rect 15764 8430 15792 11562
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15856 3233 15884 16623
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15948 10946 15976 14894
rect 16212 14748 16264 14754
rect 16212 14690 16264 14696
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 15936 10940 15988 10946
rect 15936 10882 15988 10888
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 15948 6186 15976 10746
rect 16040 6866 16068 14418
rect 16120 12912 16172 12918
rect 16120 12854 16172 12860
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 16132 3505 16160 12854
rect 16224 9858 16252 14690
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 16212 9852 16264 9858
rect 16212 9794 16264 9800
rect 16316 4321 16344 10474
rect 16302 4312 16358 4321
rect 16302 4247 16358 4256
rect 16118 3496 16174 3505
rect 16118 3431 16174 3440
rect 15842 3224 15898 3233
rect 15842 3159 15898 3168
rect 15290 2000 15346 2009
rect 15290 1935 15346 1944
rect 12346 1456 12402 1465
rect 12346 1391 12402 1400
rect 16408 921 16436 12310
rect 16500 9586 16528 12378
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 11702 912 11758 921
rect 11702 847 11758 856
rect 16394 912 16450 921
rect 16394 847 16450 856
rect 11716 513 11744 847
rect 16500 785 16528 8570
rect 16592 2689 16620 11834
rect 16684 11422 16712 16895
rect 16946 16688 17002 16697
rect 16946 16623 17002 16632
rect 16854 15600 16910 15609
rect 16854 15535 16910 15544
rect 16762 14954 16818 14963
rect 16762 14889 16818 14898
rect 16672 11416 16724 11422
rect 16672 11358 16724 11364
rect 16776 10418 16804 14889
rect 16684 10390 16804 10418
rect 16684 4049 16712 10390
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16670 4040 16726 4049
rect 16670 3975 16726 3984
rect 16578 2680 16634 2689
rect 16578 2615 16634 2624
rect 16486 776 16542 785
rect 16486 711 16542 720
rect 11702 504 11758 513
rect 11702 439 11758 448
rect 16776 377 16804 10202
rect 16868 9790 16896 15535
rect 16856 9784 16908 9790
rect 16856 9726 16908 9732
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16868 6848 16896 9522
rect 16960 7002 16988 16623
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 16868 6820 17080 6848
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16868 649 16896 6190
rect 17052 4185 17080 6820
rect 17038 4176 17094 4185
rect 17038 4111 17094 4120
rect 16854 640 16910 649
rect 16854 575 16910 584
rect 16762 368 16818 377
rect 16762 303 16818 312
rect 6918 232 6974 241
rect 6918 167 6974 176
rect 11150 232 11206 241
rect 11150 167 11206 176
<< via2 >>
rect 2410 16904 2466 16960
rect 1214 15544 1270 15600
rect 110 14864 166 14920
rect 18 12824 74 12880
rect 18 5616 74 5672
rect 386 14048 442 14104
rect 294 13776 350 13832
rect 202 11056 258 11112
rect 110 1556 166 1592
rect 110 1536 112 1556
rect 112 1536 164 1556
rect 164 1536 166 1556
rect 202 1400 258 1456
rect 662 14456 718 14512
rect 570 14320 626 14376
rect 478 1536 534 1592
rect 754 13232 810 13288
rect 938 12416 994 12472
rect 1122 8336 1178 8392
rect 1766 15444 1768 15464
rect 1768 15444 1820 15464
rect 1820 15444 1822 15464
rect 1766 15408 1822 15444
rect 2572 15802 2628 15804
rect 2652 15802 2708 15804
rect 2732 15802 2788 15804
rect 2812 15802 2868 15804
rect 2572 15750 2618 15802
rect 2618 15750 2628 15802
rect 2652 15750 2682 15802
rect 2682 15750 2694 15802
rect 2694 15750 2708 15802
rect 2732 15750 2746 15802
rect 2746 15750 2758 15802
rect 2758 15750 2788 15802
rect 2812 15750 2822 15802
rect 2822 15750 2868 15802
rect 2572 15748 2628 15750
rect 2652 15748 2708 15750
rect 2732 15748 2788 15750
rect 2812 15748 2868 15750
rect 1582 12416 1638 12472
rect 1490 11600 1546 11656
rect 3054 15308 3056 15328
rect 3056 15308 3108 15328
rect 3108 15308 3110 15328
rect 3054 15272 3110 15308
rect 2778 14884 2834 14920
rect 2778 14864 2780 14884
rect 2780 14864 2832 14884
rect 2832 14864 2834 14884
rect 2572 14714 2628 14716
rect 2652 14714 2708 14716
rect 2732 14714 2788 14716
rect 2812 14714 2868 14716
rect 2572 14662 2618 14714
rect 2618 14662 2628 14714
rect 2652 14662 2682 14714
rect 2682 14662 2694 14714
rect 2694 14662 2708 14714
rect 2732 14662 2746 14714
rect 2746 14662 2758 14714
rect 2758 14662 2788 14714
rect 2812 14662 2822 14714
rect 2822 14662 2868 14714
rect 2572 14660 2628 14662
rect 2652 14660 2708 14662
rect 2732 14660 2788 14662
rect 2812 14660 2868 14662
rect 2778 14048 2834 14104
rect 2594 13912 2650 13968
rect 3054 13776 3110 13832
rect 2572 13626 2628 13628
rect 2652 13626 2708 13628
rect 2732 13626 2788 13628
rect 2812 13626 2868 13628
rect 2572 13574 2618 13626
rect 2618 13574 2628 13626
rect 2652 13574 2682 13626
rect 2682 13574 2694 13626
rect 2694 13574 2708 13626
rect 2732 13574 2746 13626
rect 2746 13574 2758 13626
rect 2758 13574 2788 13626
rect 2812 13574 2822 13626
rect 2822 13574 2868 13626
rect 2572 13572 2628 13574
rect 2652 13572 2708 13574
rect 2732 13572 2788 13574
rect 2812 13572 2868 13574
rect 2594 12724 2596 12744
rect 2596 12724 2648 12744
rect 2648 12724 2650 12744
rect 2594 12688 2650 12724
rect 2572 12538 2628 12540
rect 2652 12538 2708 12540
rect 2732 12538 2788 12540
rect 2812 12538 2868 12540
rect 2572 12486 2618 12538
rect 2618 12486 2628 12538
rect 2652 12486 2682 12538
rect 2682 12486 2694 12538
rect 2694 12486 2708 12538
rect 2732 12486 2746 12538
rect 2746 12486 2758 12538
rect 2758 12486 2788 12538
rect 2812 12486 2822 12538
rect 2822 12486 2868 12538
rect 2572 12484 2628 12486
rect 2652 12484 2708 12486
rect 2732 12484 2788 12486
rect 2812 12484 2868 12486
rect 2042 10104 2098 10160
rect 3238 15544 3294 15600
rect 4066 16632 4122 16688
rect 6366 16768 6422 16824
rect 4066 15272 4122 15328
rect 3572 15258 3628 15260
rect 3652 15258 3708 15260
rect 3732 15258 3788 15260
rect 3812 15258 3868 15260
rect 3572 15206 3618 15258
rect 3618 15206 3628 15258
rect 3652 15206 3682 15258
rect 3682 15206 3694 15258
rect 3694 15206 3708 15258
rect 3732 15206 3746 15258
rect 3746 15206 3758 15258
rect 3758 15206 3788 15258
rect 3812 15206 3822 15258
rect 3822 15206 3868 15258
rect 3572 15204 3628 15206
rect 3652 15204 3708 15206
rect 3732 15204 3788 15206
rect 3812 15204 3868 15206
rect 3606 14320 3662 14376
rect 3572 14170 3628 14172
rect 3652 14170 3708 14172
rect 3732 14170 3788 14172
rect 3812 14170 3868 14172
rect 3572 14118 3618 14170
rect 3618 14118 3628 14170
rect 3652 14118 3682 14170
rect 3682 14118 3694 14170
rect 3694 14118 3708 14170
rect 3732 14118 3746 14170
rect 3746 14118 3758 14170
rect 3758 14118 3788 14170
rect 3812 14118 3822 14170
rect 3822 14118 3868 14170
rect 3572 14116 3628 14118
rect 3652 14116 3708 14118
rect 3732 14116 3788 14118
rect 3812 14116 3868 14118
rect 3330 12860 3332 12880
rect 3332 12860 3384 12880
rect 3384 12860 3386 12880
rect 3330 12824 3386 12860
rect 3330 12552 3386 12608
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2502 10548 2504 10568
rect 2504 10548 2556 10568
rect 2556 10548 2558 10568
rect 2502 10512 2558 10548
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 1950 5752 2006 5808
rect 3054 10240 3110 10296
rect 3146 9968 3202 10024
rect 3514 13368 3570 13424
rect 3572 13082 3628 13084
rect 3652 13082 3708 13084
rect 3732 13082 3788 13084
rect 3812 13082 3868 13084
rect 3572 13030 3618 13082
rect 3618 13030 3628 13082
rect 3652 13030 3682 13082
rect 3682 13030 3694 13082
rect 3694 13030 3708 13082
rect 3732 13030 3746 13082
rect 3746 13030 3758 13082
rect 3758 13030 3788 13082
rect 3812 13030 3822 13082
rect 3822 13030 3868 13082
rect 3572 13028 3628 13030
rect 3652 13028 3708 13030
rect 3732 13028 3788 13030
rect 3812 13028 3868 13030
rect 3572 11994 3628 11996
rect 3652 11994 3708 11996
rect 3732 11994 3788 11996
rect 3812 11994 3868 11996
rect 3572 11942 3618 11994
rect 3618 11942 3628 11994
rect 3652 11942 3682 11994
rect 3682 11942 3694 11994
rect 3694 11942 3708 11994
rect 3732 11942 3746 11994
rect 3746 11942 3758 11994
rect 3758 11942 3788 11994
rect 3812 11942 3822 11994
rect 3822 11942 3868 11994
rect 3572 11940 3628 11942
rect 3652 11940 3708 11942
rect 3732 11940 3788 11942
rect 3812 11940 3868 11942
rect 3422 11192 3478 11248
rect 3572 10906 3628 10908
rect 3652 10906 3708 10908
rect 3732 10906 3788 10908
rect 3812 10906 3868 10908
rect 3572 10854 3618 10906
rect 3618 10854 3628 10906
rect 3652 10854 3682 10906
rect 3682 10854 3694 10906
rect 3694 10854 3708 10906
rect 3732 10854 3746 10906
rect 3746 10854 3758 10906
rect 3758 10854 3788 10906
rect 3812 10854 3822 10906
rect 3822 10854 3868 10906
rect 3572 10852 3628 10854
rect 3652 10852 3708 10854
rect 3732 10852 3788 10854
rect 3812 10852 3868 10854
rect 2686 9460 2688 9480
rect 2688 9460 2740 9480
rect 2740 9460 2742 9480
rect 2134 5344 2190 5400
rect 1858 4528 1914 4584
rect 2686 9424 2742 9460
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2778 8372 2780 8392
rect 2780 8372 2832 8392
rect 2832 8372 2834 8392
rect 2778 8336 2834 8372
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2318 7792 2374 7848
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 3054 9152 3110 9208
rect 2410 6296 2466 6352
rect 3054 6024 3110 6080
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 2502 5616 2558 5672
rect 2410 4120 2466 4176
rect 2410 3984 2466 4040
rect 2686 3984 2742 4040
rect 2594 3712 2650 3768
rect 2686 3576 2742 3632
rect 3238 9696 3294 9752
rect 3238 8200 3294 8256
rect 3238 7248 3294 7304
rect 3146 3032 3202 3088
rect 2410 2488 2466 2544
rect 2410 1672 2466 1728
rect 1858 1536 1914 1592
rect 2318 1536 2374 1592
rect 2778 1400 2834 1456
rect 2962 1420 3018 1456
rect 2962 1400 2964 1420
rect 2964 1400 3016 1420
rect 3016 1400 3018 1420
rect 1122 1264 1178 1320
rect 3572 9818 3628 9820
rect 3652 9818 3708 9820
rect 3732 9818 3788 9820
rect 3812 9818 3868 9820
rect 3572 9766 3618 9818
rect 3618 9766 3628 9818
rect 3652 9766 3682 9818
rect 3682 9766 3694 9818
rect 3694 9766 3708 9818
rect 3732 9766 3746 9818
rect 3746 9766 3758 9818
rect 3758 9766 3788 9818
rect 3812 9766 3822 9818
rect 3822 9766 3868 9818
rect 3572 9764 3628 9766
rect 3652 9764 3708 9766
rect 3732 9764 3788 9766
rect 3812 9764 3868 9766
rect 4250 13232 4306 13288
rect 4710 15564 4766 15600
rect 4710 15544 4712 15564
rect 4712 15544 4764 15564
rect 4764 15544 4766 15564
rect 4342 12824 4398 12880
rect 4066 12044 4068 12064
rect 4068 12044 4120 12064
rect 4120 12044 4122 12064
rect 4066 12008 4122 12044
rect 4158 11636 4160 11656
rect 4160 11636 4212 11656
rect 4212 11636 4214 11656
rect 4158 11600 4214 11636
rect 4158 11076 4214 11112
rect 4158 11056 4160 11076
rect 4160 11056 4212 11076
rect 4212 11056 4214 11076
rect 4802 14476 4858 14512
rect 4802 14456 4804 14476
rect 4804 14456 4856 14476
rect 4856 14456 4858 14476
rect 4894 13812 4896 13832
rect 4896 13812 4948 13832
rect 4948 13812 4950 13832
rect 4894 13776 4950 13812
rect 5262 15408 5318 15464
rect 5446 14456 5502 14512
rect 4434 9968 4490 10024
rect 3572 8730 3628 8732
rect 3652 8730 3708 8732
rect 3732 8730 3788 8732
rect 3812 8730 3868 8732
rect 3572 8678 3618 8730
rect 3618 8678 3628 8730
rect 3652 8678 3682 8730
rect 3682 8678 3694 8730
rect 3694 8678 3708 8730
rect 3732 8678 3746 8730
rect 3746 8678 3758 8730
rect 3758 8678 3788 8730
rect 3812 8678 3822 8730
rect 3822 8678 3868 8730
rect 3572 8676 3628 8678
rect 3652 8676 3708 8678
rect 3732 8676 3788 8678
rect 3812 8676 3868 8678
rect 3882 8336 3938 8392
rect 3572 7642 3628 7644
rect 3652 7642 3708 7644
rect 3732 7642 3788 7644
rect 3812 7642 3868 7644
rect 3572 7590 3618 7642
rect 3618 7590 3628 7642
rect 3652 7590 3682 7642
rect 3682 7590 3694 7642
rect 3694 7590 3708 7642
rect 3732 7590 3746 7642
rect 3746 7590 3758 7642
rect 3758 7590 3788 7642
rect 3812 7590 3822 7642
rect 3822 7590 3868 7642
rect 3572 7588 3628 7590
rect 3652 7588 3708 7590
rect 3732 7588 3788 7590
rect 3812 7588 3868 7590
rect 3572 6554 3628 6556
rect 3652 6554 3708 6556
rect 3732 6554 3788 6556
rect 3812 6554 3868 6556
rect 3572 6502 3618 6554
rect 3618 6502 3628 6554
rect 3652 6502 3682 6554
rect 3682 6502 3694 6554
rect 3694 6502 3708 6554
rect 3732 6502 3746 6554
rect 3746 6502 3758 6554
rect 3758 6502 3788 6554
rect 3812 6502 3822 6554
rect 3822 6502 3868 6554
rect 3572 6500 3628 6502
rect 3652 6500 3708 6502
rect 3732 6500 3788 6502
rect 3812 6500 3868 6502
rect 3422 5616 3478 5672
rect 3330 5344 3386 5400
rect 3330 3848 3386 3904
rect 3572 5466 3628 5468
rect 3652 5466 3708 5468
rect 3732 5466 3788 5468
rect 3812 5466 3868 5468
rect 3572 5414 3618 5466
rect 3618 5414 3628 5466
rect 3652 5414 3682 5466
rect 3682 5414 3694 5466
rect 3694 5414 3708 5466
rect 3732 5414 3746 5466
rect 3746 5414 3758 5466
rect 3758 5414 3788 5466
rect 3812 5414 3822 5466
rect 3822 5414 3868 5466
rect 3572 5412 3628 5414
rect 3652 5412 3708 5414
rect 3732 5412 3788 5414
rect 3812 5412 3868 5414
rect 4066 6976 4122 7032
rect 4434 9288 4490 9344
rect 4342 5616 4398 5672
rect 3514 4664 3570 4720
rect 3572 4378 3628 4380
rect 3652 4378 3708 4380
rect 3732 4378 3788 4380
rect 3812 4378 3868 4380
rect 3572 4326 3618 4378
rect 3618 4326 3628 4378
rect 3652 4326 3682 4378
rect 3682 4326 3694 4378
rect 3694 4326 3708 4378
rect 3732 4326 3746 4378
rect 3746 4326 3758 4378
rect 3758 4326 3788 4378
rect 3812 4326 3822 4378
rect 3822 4326 3868 4378
rect 3572 4324 3628 4326
rect 3652 4324 3708 4326
rect 3732 4324 3788 4326
rect 3812 4324 3868 4326
rect 4158 4392 4214 4448
rect 4066 4140 4122 4176
rect 4066 4120 4068 4140
rect 4068 4120 4120 4140
rect 4120 4120 4122 4140
rect 3572 3290 3628 3292
rect 3652 3290 3708 3292
rect 3732 3290 3788 3292
rect 3812 3290 3868 3292
rect 3572 3238 3618 3290
rect 3618 3238 3628 3290
rect 3652 3238 3682 3290
rect 3682 3238 3694 3290
rect 3694 3238 3708 3290
rect 3732 3238 3746 3290
rect 3746 3238 3758 3290
rect 3758 3238 3788 3290
rect 3812 3238 3822 3290
rect 3822 3238 3868 3290
rect 3572 3236 3628 3238
rect 3652 3236 3708 3238
rect 3732 3236 3788 3238
rect 3812 3236 3868 3238
rect 3572 2202 3628 2204
rect 3652 2202 3708 2204
rect 3732 2202 3788 2204
rect 3812 2202 3868 2204
rect 3572 2150 3618 2202
rect 3618 2150 3628 2202
rect 3652 2150 3682 2202
rect 3682 2150 3694 2202
rect 3694 2150 3708 2202
rect 3732 2150 3746 2202
rect 3746 2150 3758 2202
rect 3758 2150 3788 2202
rect 3812 2150 3822 2202
rect 3822 2150 3868 2202
rect 3572 2148 3628 2150
rect 3652 2148 3708 2150
rect 3732 2148 3788 2150
rect 3812 2148 3868 2150
rect 4066 3984 4122 4040
rect 4066 2624 4122 2680
rect 4894 12280 4950 12336
rect 4986 11056 5042 11112
rect 4894 10648 4950 10704
rect 4710 5752 4766 5808
rect 4894 5208 4950 5264
rect 4710 3052 4766 3088
rect 4710 3032 4712 3052
rect 4712 3032 4764 3052
rect 4764 3032 4766 3052
rect 4158 1536 4214 1592
rect 3606 1300 3608 1320
rect 3608 1300 3660 1320
rect 3660 1300 3662 1320
rect 3606 1264 3662 1300
rect 4066 1284 4122 1320
rect 4066 1264 4068 1284
rect 4068 1264 4120 1284
rect 4120 1264 4122 1284
rect 570 1128 626 1184
rect 3422 1128 3478 1184
rect 3572 1114 3628 1116
rect 3652 1114 3708 1116
rect 3732 1114 3788 1116
rect 3812 1114 3868 1116
rect 3572 1062 3618 1114
rect 3618 1062 3628 1114
rect 3652 1062 3682 1114
rect 3682 1062 3694 1114
rect 3694 1062 3708 1114
rect 3732 1062 3746 1114
rect 3746 1062 3758 1114
rect 3758 1062 3788 1114
rect 3812 1062 3822 1114
rect 3822 1062 3868 1114
rect 3572 1060 3628 1062
rect 3652 1060 3708 1062
rect 3732 1060 3788 1062
rect 3812 1060 3868 1062
rect 386 856 442 912
rect 5538 12552 5594 12608
rect 5170 8064 5226 8120
rect 5354 8880 5410 8936
rect 5906 13368 5962 13424
rect 16670 16904 16726 16960
rect 13358 16768 13414 16824
rect 6826 16088 6882 16144
rect 10874 16088 10930 16144
rect 7572 15802 7628 15804
rect 7652 15802 7708 15804
rect 7732 15802 7788 15804
rect 7812 15802 7868 15804
rect 7572 15750 7618 15802
rect 7618 15750 7628 15802
rect 7652 15750 7682 15802
rect 7682 15750 7694 15802
rect 7694 15750 7708 15802
rect 7732 15750 7746 15802
rect 7746 15750 7758 15802
rect 7758 15750 7788 15802
rect 7812 15750 7822 15802
rect 7822 15750 7868 15802
rect 7572 15748 7628 15750
rect 7652 15748 7708 15750
rect 7732 15748 7788 15750
rect 7812 15748 7868 15750
rect 8114 15428 8170 15464
rect 8114 15408 8116 15428
rect 8116 15408 8168 15428
rect 8168 15408 8170 15428
rect 6642 15308 6644 15328
rect 6644 15308 6696 15328
rect 6696 15308 6698 15328
rect 6642 15272 6698 15308
rect 6550 15136 6606 15192
rect 8572 15258 8628 15260
rect 8652 15258 8708 15260
rect 8732 15258 8788 15260
rect 8812 15258 8868 15260
rect 8572 15206 8618 15258
rect 8618 15206 8628 15258
rect 8652 15206 8682 15258
rect 8682 15206 8694 15258
rect 8694 15206 8708 15258
rect 8732 15206 8746 15258
rect 8746 15206 8758 15258
rect 8758 15206 8788 15258
rect 8812 15206 8822 15258
rect 8822 15206 8868 15258
rect 8572 15204 8628 15206
rect 8652 15204 8708 15206
rect 8732 15204 8788 15206
rect 8812 15204 8868 15206
rect 8390 15136 8446 15192
rect 7102 14320 7158 14376
rect 5998 12280 6054 12336
rect 5906 12164 5962 12200
rect 5906 12144 5908 12164
rect 5908 12144 5960 12164
rect 5960 12144 5962 12164
rect 5722 10240 5778 10296
rect 5630 10104 5686 10160
rect 5630 8472 5686 8528
rect 5538 7792 5594 7848
rect 5170 6840 5226 6896
rect 5538 7112 5594 7168
rect 5814 10104 5870 10160
rect 5998 9696 6054 9752
rect 5814 9560 5870 9616
rect 5814 8744 5870 8800
rect 5906 8336 5962 8392
rect 5354 5888 5410 5944
rect 5354 4800 5410 4856
rect 5722 6704 5778 6760
rect 5722 4528 5778 4584
rect 5446 3712 5502 3768
rect 5630 3576 5686 3632
rect 5078 3304 5134 3360
rect 5354 3052 5410 3088
rect 5354 3032 5356 3052
rect 5356 3032 5408 3052
rect 5408 3032 5410 3052
rect 5630 2524 5632 2544
rect 5632 2524 5684 2544
rect 5684 2524 5686 2544
rect 5630 2488 5686 2524
rect 5630 2352 5686 2408
rect 5446 1536 5502 1592
rect 7572 14714 7628 14716
rect 7652 14714 7708 14716
rect 7732 14714 7788 14716
rect 7812 14714 7868 14716
rect 7572 14662 7618 14714
rect 7618 14662 7628 14714
rect 7652 14662 7682 14714
rect 7682 14662 7694 14714
rect 7694 14662 7708 14714
rect 7732 14662 7746 14714
rect 7746 14662 7758 14714
rect 7758 14662 7788 14714
rect 7812 14662 7822 14714
rect 7822 14662 7868 14714
rect 7572 14660 7628 14662
rect 7652 14660 7708 14662
rect 7732 14660 7788 14662
rect 7812 14660 7868 14662
rect 8942 14864 8998 14920
rect 6918 12008 6974 12064
rect 7010 11056 7066 11112
rect 6366 6976 6422 7032
rect 6274 6840 6330 6896
rect 6182 5888 6238 5944
rect 6182 5616 6238 5672
rect 5998 4700 6000 4720
rect 6000 4700 6052 4720
rect 6052 4700 6054 4720
rect 5998 4664 6054 4700
rect 5998 4528 6054 4584
rect 7010 9832 7066 9888
rect 7010 9288 7066 9344
rect 7194 11076 7250 11112
rect 7194 11056 7196 11076
rect 7196 11056 7248 11076
rect 7248 11056 7250 11076
rect 7102 8200 7158 8256
rect 6642 6160 6698 6216
rect 6550 5752 6606 5808
rect 7102 7112 7158 7168
rect 6182 3884 6184 3904
rect 6184 3884 6236 3904
rect 6236 3884 6238 3904
rect 6182 3848 6238 3884
rect 7572 13626 7628 13628
rect 7652 13626 7708 13628
rect 7732 13626 7788 13628
rect 7812 13626 7868 13628
rect 7572 13574 7618 13626
rect 7618 13574 7628 13626
rect 7652 13574 7682 13626
rect 7682 13574 7694 13626
rect 7694 13574 7708 13626
rect 7732 13574 7746 13626
rect 7746 13574 7758 13626
rect 7758 13574 7788 13626
rect 7812 13574 7822 13626
rect 7822 13574 7868 13626
rect 7572 13572 7628 13574
rect 7652 13572 7708 13574
rect 7732 13572 7788 13574
rect 7812 13572 7868 13574
rect 7572 12538 7628 12540
rect 7652 12538 7708 12540
rect 7732 12538 7788 12540
rect 7812 12538 7868 12540
rect 7572 12486 7618 12538
rect 7618 12486 7628 12538
rect 7652 12486 7682 12538
rect 7682 12486 7694 12538
rect 7694 12486 7708 12538
rect 7732 12486 7746 12538
rect 7746 12486 7758 12538
rect 7758 12486 7788 12538
rect 7812 12486 7822 12538
rect 7822 12486 7868 12538
rect 7572 12484 7628 12486
rect 7652 12484 7708 12486
rect 7732 12484 7788 12486
rect 7812 12484 7868 12486
rect 7572 11450 7628 11452
rect 7652 11450 7708 11452
rect 7732 11450 7788 11452
rect 7812 11450 7868 11452
rect 7572 11398 7618 11450
rect 7618 11398 7628 11450
rect 7652 11398 7682 11450
rect 7682 11398 7694 11450
rect 7694 11398 7708 11450
rect 7732 11398 7746 11450
rect 7746 11398 7758 11450
rect 7758 11398 7788 11450
rect 7812 11398 7822 11450
rect 7822 11398 7868 11450
rect 7572 11396 7628 11398
rect 7652 11396 7708 11398
rect 7732 11396 7788 11398
rect 7812 11396 7868 11398
rect 8022 13912 8078 13968
rect 8114 13096 8170 13152
rect 8206 12824 8262 12880
rect 7572 10362 7628 10364
rect 7652 10362 7708 10364
rect 7732 10362 7788 10364
rect 7812 10362 7868 10364
rect 7572 10310 7618 10362
rect 7618 10310 7628 10362
rect 7652 10310 7682 10362
rect 7682 10310 7694 10362
rect 7694 10310 7708 10362
rect 7732 10310 7746 10362
rect 7746 10310 7758 10362
rect 7758 10310 7788 10362
rect 7812 10310 7822 10362
rect 7822 10310 7868 10362
rect 7572 10308 7628 10310
rect 7652 10308 7708 10310
rect 7732 10308 7788 10310
rect 7812 10308 7868 10310
rect 8022 9968 8078 10024
rect 7194 6024 7250 6080
rect 7194 5072 7250 5128
rect 5998 3440 6054 3496
rect 6090 2488 6146 2544
rect 6274 1944 6330 2000
rect 6550 1672 6606 1728
rect 4710 856 4766 912
rect 4894 856 4950 912
rect 4342 720 4398 776
rect 7010 3576 7066 3632
rect 7572 9274 7628 9276
rect 7652 9274 7708 9276
rect 7732 9274 7788 9276
rect 7812 9274 7868 9276
rect 7572 9222 7618 9274
rect 7618 9222 7628 9274
rect 7652 9222 7682 9274
rect 7682 9222 7694 9274
rect 7694 9222 7708 9274
rect 7732 9222 7746 9274
rect 7746 9222 7758 9274
rect 7758 9222 7788 9274
rect 7812 9222 7822 9274
rect 7822 9222 7868 9274
rect 7572 9220 7628 9222
rect 7652 9220 7708 9222
rect 7732 9220 7788 9222
rect 7812 9220 7868 9222
rect 8022 9152 8078 9208
rect 8022 8744 8078 8800
rect 7572 8186 7628 8188
rect 7652 8186 7708 8188
rect 7732 8186 7788 8188
rect 7812 8186 7868 8188
rect 7572 8134 7618 8186
rect 7618 8134 7628 8186
rect 7652 8134 7682 8186
rect 7682 8134 7694 8186
rect 7694 8134 7708 8186
rect 7732 8134 7746 8186
rect 7746 8134 7758 8186
rect 7758 8134 7788 8186
rect 7812 8134 7822 8186
rect 7822 8134 7868 8186
rect 7572 8132 7628 8134
rect 7652 8132 7708 8134
rect 7732 8132 7788 8134
rect 7812 8132 7868 8134
rect 8572 14170 8628 14172
rect 8652 14170 8708 14172
rect 8732 14170 8788 14172
rect 8812 14170 8868 14172
rect 8572 14118 8618 14170
rect 8618 14118 8628 14170
rect 8652 14118 8682 14170
rect 8682 14118 8694 14170
rect 8694 14118 8708 14170
rect 8732 14118 8746 14170
rect 8746 14118 8758 14170
rect 8758 14118 8788 14170
rect 8812 14118 8822 14170
rect 8822 14118 8868 14170
rect 8572 14116 8628 14118
rect 8652 14116 8708 14118
rect 8732 14116 8788 14118
rect 8812 14116 8868 14118
rect 8942 13932 8998 13968
rect 8942 13912 8944 13932
rect 8944 13912 8996 13932
rect 8996 13912 8998 13932
rect 8572 13082 8628 13084
rect 8652 13082 8708 13084
rect 8732 13082 8788 13084
rect 8812 13082 8868 13084
rect 8572 13030 8618 13082
rect 8618 13030 8628 13082
rect 8652 13030 8682 13082
rect 8682 13030 8694 13082
rect 8694 13030 8708 13082
rect 8732 13030 8746 13082
rect 8746 13030 8758 13082
rect 8758 13030 8788 13082
rect 8812 13030 8822 13082
rect 8822 13030 8868 13082
rect 8572 13028 8628 13030
rect 8652 13028 8708 13030
rect 8732 13028 8788 13030
rect 8812 13028 8868 13030
rect 8942 12280 8998 12336
rect 8572 11994 8628 11996
rect 8652 11994 8708 11996
rect 8732 11994 8788 11996
rect 8812 11994 8868 11996
rect 8572 11942 8618 11994
rect 8618 11942 8628 11994
rect 8652 11942 8682 11994
rect 8682 11942 8694 11994
rect 8694 11942 8708 11994
rect 8732 11942 8746 11994
rect 8746 11942 8758 11994
rect 8758 11942 8788 11994
rect 8812 11942 8822 11994
rect 8822 11942 8868 11994
rect 8572 11940 8628 11942
rect 8652 11940 8708 11942
rect 8732 11940 8788 11942
rect 8812 11940 8868 11942
rect 9126 15308 9128 15328
rect 9128 15308 9180 15328
rect 9180 15308 9182 15328
rect 9126 15272 9182 15308
rect 10690 14864 10746 14920
rect 9310 14048 9366 14104
rect 8850 11772 8852 11792
rect 8852 11772 8904 11792
rect 8904 11772 8906 11792
rect 8850 11736 8906 11772
rect 8758 11328 8814 11384
rect 8572 10906 8628 10908
rect 8652 10906 8708 10908
rect 8732 10906 8788 10908
rect 8812 10906 8868 10908
rect 8572 10854 8618 10906
rect 8618 10854 8628 10906
rect 8652 10854 8682 10906
rect 8682 10854 8694 10906
rect 8694 10854 8708 10906
rect 8732 10854 8746 10906
rect 8746 10854 8758 10906
rect 8758 10854 8788 10906
rect 8812 10854 8822 10906
rect 8822 10854 8868 10906
rect 8572 10852 8628 10854
rect 8652 10852 8708 10854
rect 8732 10852 8788 10854
rect 8812 10852 8868 10854
rect 8206 9832 8262 9888
rect 8298 9696 8354 9752
rect 8206 8372 8208 8392
rect 8208 8372 8260 8392
rect 8260 8372 8262 8392
rect 8206 8336 8262 8372
rect 7572 7098 7628 7100
rect 7652 7098 7708 7100
rect 7732 7098 7788 7100
rect 7812 7098 7868 7100
rect 7572 7046 7618 7098
rect 7618 7046 7628 7098
rect 7652 7046 7682 7098
rect 7682 7046 7694 7098
rect 7694 7046 7708 7098
rect 7732 7046 7746 7098
rect 7746 7046 7758 7098
rect 7758 7046 7788 7098
rect 7812 7046 7822 7098
rect 7822 7046 7868 7098
rect 7572 7044 7628 7046
rect 7652 7044 7708 7046
rect 7732 7044 7788 7046
rect 7812 7044 7868 7046
rect 7286 4800 7342 4856
rect 7572 6010 7628 6012
rect 7652 6010 7708 6012
rect 7732 6010 7788 6012
rect 7812 6010 7868 6012
rect 7572 5958 7618 6010
rect 7618 5958 7628 6010
rect 7652 5958 7682 6010
rect 7682 5958 7694 6010
rect 7694 5958 7708 6010
rect 7732 5958 7746 6010
rect 7746 5958 7758 6010
rect 7758 5958 7788 6010
rect 7812 5958 7822 6010
rect 7822 5958 7868 6010
rect 7572 5956 7628 5958
rect 7652 5956 7708 5958
rect 7732 5956 7788 5958
rect 7812 5956 7868 5958
rect 7572 4922 7628 4924
rect 7652 4922 7708 4924
rect 7732 4922 7788 4924
rect 7812 4922 7868 4924
rect 7572 4870 7618 4922
rect 7618 4870 7628 4922
rect 7652 4870 7682 4922
rect 7682 4870 7694 4922
rect 7694 4870 7708 4922
rect 7732 4870 7746 4922
rect 7746 4870 7758 4922
rect 7758 4870 7788 4922
rect 7812 4870 7822 4922
rect 7822 4870 7868 4922
rect 7572 4868 7628 4870
rect 7652 4868 7708 4870
rect 7732 4868 7788 4870
rect 7812 4868 7868 4870
rect 7572 3834 7628 3836
rect 7652 3834 7708 3836
rect 7732 3834 7788 3836
rect 7812 3834 7868 3836
rect 7572 3782 7618 3834
rect 7618 3782 7628 3834
rect 7652 3782 7682 3834
rect 7682 3782 7694 3834
rect 7694 3782 7708 3834
rect 7732 3782 7746 3834
rect 7746 3782 7758 3834
rect 7758 3782 7788 3834
rect 7812 3782 7822 3834
rect 7822 3782 7868 3834
rect 7572 3780 7628 3782
rect 7652 3780 7708 3782
rect 7732 3780 7788 3782
rect 7812 3780 7868 3782
rect 8206 6024 8262 6080
rect 8390 6840 8446 6896
rect 8206 4428 8208 4448
rect 8208 4428 8260 4448
rect 8260 4428 8262 4448
rect 8206 4392 8262 4428
rect 8206 3712 8262 3768
rect 9310 12552 9366 12608
rect 8572 9818 8628 9820
rect 8652 9818 8708 9820
rect 8732 9818 8788 9820
rect 8812 9818 8868 9820
rect 8572 9766 8618 9818
rect 8618 9766 8628 9818
rect 8652 9766 8682 9818
rect 8682 9766 8694 9818
rect 8694 9766 8708 9818
rect 8732 9766 8746 9818
rect 8746 9766 8758 9818
rect 8758 9766 8788 9818
rect 8812 9766 8822 9818
rect 8822 9766 8868 9818
rect 8572 9764 8628 9766
rect 8652 9764 8708 9766
rect 8732 9764 8788 9766
rect 8812 9764 8868 9766
rect 8942 9560 8998 9616
rect 9218 10648 9274 10704
rect 9126 9868 9128 9888
rect 9128 9868 9180 9888
rect 9180 9868 9182 9888
rect 9126 9832 9182 9868
rect 8942 8880 8998 8936
rect 8572 8730 8628 8732
rect 8652 8730 8708 8732
rect 8732 8730 8788 8732
rect 8812 8730 8868 8732
rect 8572 8678 8618 8730
rect 8618 8678 8628 8730
rect 8652 8678 8682 8730
rect 8682 8678 8694 8730
rect 8694 8678 8708 8730
rect 8732 8678 8746 8730
rect 8746 8678 8758 8730
rect 8758 8678 8788 8730
rect 8812 8678 8822 8730
rect 8822 8678 8868 8730
rect 8572 8676 8628 8678
rect 8652 8676 8708 8678
rect 8732 8676 8788 8678
rect 8812 8676 8868 8678
rect 8572 7642 8628 7644
rect 8652 7642 8708 7644
rect 8732 7642 8788 7644
rect 8812 7642 8868 7644
rect 8572 7590 8618 7642
rect 8618 7590 8628 7642
rect 8652 7590 8682 7642
rect 8682 7590 8694 7642
rect 8694 7590 8708 7642
rect 8732 7590 8746 7642
rect 8746 7590 8758 7642
rect 8758 7590 8788 7642
rect 8812 7590 8822 7642
rect 8822 7590 8868 7642
rect 8572 7588 8628 7590
rect 8652 7588 8708 7590
rect 8732 7588 8788 7590
rect 8812 7588 8868 7590
rect 8572 6554 8628 6556
rect 8652 6554 8708 6556
rect 8732 6554 8788 6556
rect 8812 6554 8868 6556
rect 8572 6502 8618 6554
rect 8618 6502 8628 6554
rect 8652 6502 8682 6554
rect 8682 6502 8694 6554
rect 8694 6502 8708 6554
rect 8732 6502 8746 6554
rect 8746 6502 8758 6554
rect 8758 6502 8788 6554
rect 8812 6502 8822 6554
rect 8822 6502 8868 6554
rect 8572 6500 8628 6502
rect 8652 6500 8708 6502
rect 8732 6500 8788 6502
rect 8812 6500 8868 6502
rect 8850 5616 8906 5672
rect 8572 5466 8628 5468
rect 8652 5466 8708 5468
rect 8732 5466 8788 5468
rect 8812 5466 8868 5468
rect 8572 5414 8618 5466
rect 8618 5414 8628 5466
rect 8652 5414 8682 5466
rect 8682 5414 8694 5466
rect 8694 5414 8708 5466
rect 8732 5414 8746 5466
rect 8746 5414 8758 5466
rect 8758 5414 8788 5466
rect 8812 5414 8822 5466
rect 8822 5414 8868 5466
rect 8572 5412 8628 5414
rect 8652 5412 8708 5414
rect 8732 5412 8788 5414
rect 8812 5412 8868 5414
rect 8574 4936 8630 4992
rect 8572 4378 8628 4380
rect 8652 4378 8708 4380
rect 8732 4378 8788 4380
rect 8812 4378 8868 4380
rect 8572 4326 8618 4378
rect 8618 4326 8628 4378
rect 8652 4326 8682 4378
rect 8682 4326 8694 4378
rect 8694 4326 8708 4378
rect 8732 4326 8746 4378
rect 8746 4326 8758 4378
rect 8758 4326 8788 4378
rect 8812 4326 8822 4378
rect 8822 4326 8868 4378
rect 8572 4324 8628 4326
rect 8652 4324 8708 4326
rect 8732 4324 8788 4326
rect 8812 4324 8868 4326
rect 9126 6160 9182 6216
rect 10322 14340 10378 14376
rect 10322 14320 10324 14340
rect 10324 14320 10376 14340
rect 10376 14320 10378 14340
rect 9678 10784 9734 10840
rect 9494 10512 9550 10568
rect 8390 3340 8392 3360
rect 8392 3340 8444 3360
rect 8444 3340 8446 3360
rect 6826 1400 6882 1456
rect 7572 2746 7628 2748
rect 7652 2746 7708 2748
rect 7732 2746 7788 2748
rect 7812 2746 7868 2748
rect 7572 2694 7618 2746
rect 7618 2694 7628 2746
rect 7652 2694 7682 2746
rect 7682 2694 7694 2746
rect 7694 2694 7708 2746
rect 7732 2694 7746 2746
rect 7746 2694 7758 2746
rect 7758 2694 7788 2746
rect 7812 2694 7822 2746
rect 7822 2694 7868 2746
rect 7572 2692 7628 2694
rect 7652 2692 7708 2694
rect 7732 2692 7788 2694
rect 7812 2692 7868 2694
rect 8022 2760 8078 2816
rect 8022 2624 8078 2680
rect 8390 3304 8446 3340
rect 8572 3290 8628 3292
rect 8652 3290 8708 3292
rect 8732 3290 8788 3292
rect 8812 3290 8868 3292
rect 8572 3238 8618 3290
rect 8618 3238 8628 3290
rect 8652 3238 8682 3290
rect 8682 3238 8694 3290
rect 8694 3238 8708 3290
rect 8732 3238 8746 3290
rect 8746 3238 8758 3290
rect 8758 3238 8788 3290
rect 8812 3238 8822 3290
rect 8822 3238 8868 3290
rect 8572 3236 8628 3238
rect 8652 3236 8708 3238
rect 8732 3236 8788 3238
rect 8812 3236 8868 3238
rect 9218 5072 9274 5128
rect 9218 3884 9220 3904
rect 9220 3884 9272 3904
rect 9272 3884 9274 3904
rect 9218 3848 9274 3884
rect 9218 3188 9274 3224
rect 9218 3168 9220 3188
rect 9220 3168 9272 3188
rect 9272 3168 9274 3188
rect 8482 2488 8538 2544
rect 8572 2202 8628 2204
rect 8652 2202 8708 2204
rect 8732 2202 8788 2204
rect 8812 2202 8868 2204
rect 8572 2150 8618 2202
rect 8618 2150 8628 2202
rect 8652 2150 8682 2202
rect 8682 2150 8694 2202
rect 8694 2150 8708 2202
rect 8732 2150 8746 2202
rect 8746 2150 8758 2202
rect 8758 2150 8788 2202
rect 8812 2150 8822 2202
rect 8822 2150 8868 2202
rect 8572 2148 8628 2150
rect 8652 2148 8708 2150
rect 8732 2148 8788 2150
rect 8812 2148 8868 2150
rect 9678 5752 9734 5808
rect 9678 4528 9734 4584
rect 9862 5480 9918 5536
rect 11886 15952 11942 16008
rect 11058 15544 11114 15600
rect 11702 15272 11758 15328
rect 11058 14592 11114 14648
rect 11058 14048 11114 14104
rect 11058 12552 11114 12608
rect 11610 12688 11666 12744
rect 11794 12824 11850 12880
rect 11794 11872 11850 11928
rect 12898 14456 12954 14512
rect 12714 12008 12770 12064
rect 11886 11736 11942 11792
rect 12530 11328 12586 11384
rect 12438 10376 12494 10432
rect 11702 9424 11758 9480
rect 10046 9152 10102 9208
rect 11794 8200 11850 8256
rect 10506 6024 10562 6080
rect 10322 5344 10378 5400
rect 8482 1844 8484 1864
rect 8484 1844 8536 1864
rect 8536 1844 8538 1864
rect 8482 1808 8538 1844
rect 10690 3440 10746 3496
rect 10690 2352 10746 2408
rect 8666 1672 8722 1728
rect 10322 1672 10378 1728
rect 7572 1658 7628 1660
rect 7652 1658 7708 1660
rect 7732 1658 7788 1660
rect 7812 1658 7868 1660
rect 7572 1606 7618 1658
rect 7618 1606 7628 1658
rect 7652 1606 7682 1658
rect 7682 1606 7694 1658
rect 7694 1606 7708 1658
rect 7732 1606 7746 1658
rect 7746 1606 7758 1658
rect 7758 1606 7788 1658
rect 7812 1606 7822 1658
rect 7822 1606 7868 1658
rect 7572 1604 7628 1606
rect 7652 1604 7708 1606
rect 7732 1604 7788 1606
rect 7812 1604 7868 1606
rect 11058 5616 11114 5672
rect 11058 5208 11114 5264
rect 11058 4392 11114 4448
rect 11058 3576 11114 3632
rect 10874 3032 10930 3088
rect 7378 1300 7380 1320
rect 7380 1300 7432 1320
rect 7432 1300 7434 1320
rect 7378 1264 7434 1300
rect 10782 1264 10838 1320
rect 8572 1114 8628 1116
rect 8652 1114 8708 1116
rect 8732 1114 8788 1116
rect 8812 1114 8868 1116
rect 8572 1062 8618 1114
rect 8618 1062 8628 1114
rect 8652 1062 8682 1114
rect 8682 1062 8694 1114
rect 8694 1062 8708 1114
rect 8732 1062 8746 1114
rect 8746 1062 8758 1114
rect 8758 1062 8788 1114
rect 8812 1062 8822 1114
rect 8822 1062 8868 1114
rect 8572 1060 8628 1062
rect 8652 1060 8708 1062
rect 8732 1060 8788 1062
rect 8812 1060 8868 1062
rect 7102 720 7158 776
rect 7286 720 7342 776
rect 6734 584 6790 640
rect 6642 448 6698 504
rect 6918 448 6974 504
rect 7102 448 7158 504
rect 4158 312 4214 368
rect 11886 6976 11942 7032
rect 11794 6704 11850 6760
rect 11242 6568 11298 6624
rect 11334 5208 11390 5264
rect 11242 3576 11298 3632
rect 12346 6160 12402 6216
rect 11886 4664 11942 4720
rect 11794 4528 11850 4584
rect 11794 1808 11850 1864
rect 12622 9968 12678 10024
rect 12530 5208 12586 5264
rect 12438 4936 12494 4992
rect 12806 11600 12862 11656
rect 12714 5480 12770 5536
rect 12622 3712 12678 3768
rect 13174 12572 13230 12608
rect 13174 12552 13176 12572
rect 13176 12552 13228 12572
rect 13228 12552 13230 12572
rect 15842 16632 15898 16688
rect 13726 15408 13782 15464
rect 13818 14748 13874 14784
rect 13818 14728 13820 14748
rect 13820 14728 13872 14748
rect 13872 14728 13874 14748
rect 13542 13912 13598 13968
rect 13726 13912 13782 13968
rect 13450 13776 13506 13832
rect 13358 12416 13414 12472
rect 13358 11056 13414 11112
rect 13082 9832 13138 9888
rect 12990 8336 13046 8392
rect 12898 6160 12954 6216
rect 13266 7384 13322 7440
rect 12990 4936 13046 4992
rect 12806 3576 12862 3632
rect 13358 6160 13414 6216
rect 13266 3848 13322 3904
rect 13174 2896 13230 2952
rect 13450 5752 13506 5808
rect 13634 13368 13690 13424
rect 13818 13116 13874 13152
rect 13818 13096 13820 13116
rect 13820 13096 13872 13116
rect 13872 13096 13874 13116
rect 13818 11092 13820 11112
rect 13820 11092 13872 11112
rect 13872 11092 13874 11112
rect 13818 11056 13874 11092
rect 13818 10784 13874 10840
rect 13726 10648 13782 10704
rect 13818 9868 13820 9888
rect 13820 9868 13872 9888
rect 13872 9868 13874 9888
rect 13818 9832 13874 9868
rect 13818 9424 13874 9480
rect 13818 9016 13874 9072
rect 13726 7792 13782 7848
rect 13542 5616 13598 5672
rect 13818 6296 13874 6352
rect 13818 5752 13874 5808
rect 13726 5072 13782 5128
rect 13818 4836 13820 4856
rect 13820 4836 13872 4856
rect 13872 4836 13874 4856
rect 13818 4800 13874 4836
rect 13726 4392 13782 4448
rect 15152 13504 15208 13560
rect 15152 12280 15208 12336
rect 15152 11464 15208 11520
rect 15152 10240 15208 10296
rect 14554 4256 14610 4312
rect 14002 3304 14058 3360
rect 14554 2760 14610 2816
rect 16302 4256 16358 4312
rect 16118 3440 16174 3496
rect 15842 3168 15898 3224
rect 15290 1944 15346 2000
rect 12346 1400 12402 1456
rect 11702 856 11758 912
rect 16394 856 16450 912
rect 16946 16632 17002 16688
rect 16854 15544 16910 15600
rect 16762 14898 16818 14954
rect 16670 3984 16726 4040
rect 16578 2624 16634 2680
rect 16486 720 16542 776
rect 11702 448 11758 504
rect 17038 4120 17094 4176
rect 16854 584 16910 640
rect 16762 312 16818 368
rect 6918 176 6974 232
rect 11150 176 11206 232
<< metal3 >>
rect 2405 16962 2471 16965
rect 16665 16962 16731 16965
rect 2405 16960 16731 16962
rect 2405 16904 2410 16960
rect 2466 16904 16670 16960
rect 16726 16904 16731 16960
rect 2405 16902 16731 16904
rect 2405 16899 2471 16902
rect 16665 16899 16731 16902
rect 6361 16826 6427 16829
rect 13353 16826 13419 16829
rect 6361 16824 13419 16826
rect 6361 16768 6366 16824
rect 6422 16768 13358 16824
rect 13414 16768 13419 16824
rect 6361 16766 13419 16768
rect 6361 16763 6427 16766
rect 13353 16763 13419 16766
rect 4061 16690 4127 16693
rect 15837 16690 15903 16693
rect 4061 16688 15903 16690
rect 4061 16632 4066 16688
rect 4122 16632 15842 16688
rect 15898 16632 15903 16688
rect 4061 16630 15903 16632
rect 4061 16627 4127 16630
rect 15837 16627 15903 16630
rect 16941 16690 17007 16693
rect 16941 16688 17050 16690
rect 16941 16632 16946 16688
rect 17002 16632 17050 16688
rect 16941 16627 17050 16632
rect 16990 16448 17050 16627
rect 14000 16328 34000 16448
rect 6821 16146 6887 16149
rect 10869 16146 10935 16149
rect 6821 16144 10935 16146
rect 6821 16088 6826 16144
rect 6882 16088 10874 16144
rect 10930 16088 10935 16144
rect 6821 16086 10935 16088
rect 6821 16083 6887 16086
rect 10869 16083 10935 16086
rect 11881 16010 11947 16013
rect 14000 16010 34000 16040
rect 11881 16008 34000 16010
rect 11881 15952 11886 16008
rect 11942 15952 34000 16008
rect 11881 15950 34000 15952
rect 11881 15947 11947 15950
rect 14000 15920 34000 15950
rect 2562 15808 2878 15809
rect 2562 15744 2568 15808
rect 2632 15744 2648 15808
rect 2712 15744 2728 15808
rect 2792 15744 2808 15808
rect 2872 15744 2878 15808
rect 2562 15743 2878 15744
rect 7562 15808 7878 15809
rect 7562 15744 7568 15808
rect 7632 15744 7648 15808
rect 7712 15744 7728 15808
rect 7792 15744 7808 15808
rect 7872 15744 7878 15808
rect 7562 15743 7878 15744
rect 1209 15602 1275 15605
rect 3233 15602 3299 15605
rect 1209 15600 3299 15602
rect 1209 15544 1214 15600
rect 1270 15544 3238 15600
rect 3294 15544 3299 15600
rect 1209 15542 3299 15544
rect 1209 15539 1275 15542
rect 3233 15539 3299 15542
rect 4705 15602 4771 15605
rect 11053 15602 11119 15605
rect 4705 15600 11119 15602
rect 4705 15544 4710 15600
rect 4766 15544 11058 15600
rect 11114 15544 11119 15600
rect 4705 15542 11119 15544
rect 4705 15539 4771 15542
rect 11053 15539 11119 15542
rect 14000 15600 34000 15632
rect 14000 15544 16854 15600
rect 16910 15544 34000 15600
rect 14000 15512 34000 15544
rect 1761 15466 1827 15469
rect 5257 15466 5323 15469
rect 1761 15464 5323 15466
rect 1761 15408 1766 15464
rect 1822 15408 5262 15464
rect 5318 15408 5323 15464
rect 1761 15406 5323 15408
rect 1761 15403 1827 15406
rect 5257 15403 5323 15406
rect 8109 15466 8175 15469
rect 13721 15466 13787 15469
rect 8109 15464 13787 15466
rect 8109 15408 8114 15464
rect 8170 15408 13726 15464
rect 13782 15408 13787 15464
rect 8109 15406 13787 15408
rect 8109 15403 8175 15406
rect 13721 15403 13787 15406
rect 974 15268 980 15332
rect 1044 15330 1050 15332
rect 3049 15330 3115 15333
rect 1044 15328 3115 15330
rect 1044 15272 3054 15328
rect 3110 15272 3115 15328
rect 1044 15270 3115 15272
rect 1044 15268 1050 15270
rect 3049 15267 3115 15270
rect 4061 15330 4127 15333
rect 6637 15330 6703 15333
rect 4061 15328 6703 15330
rect 4061 15272 4066 15328
rect 4122 15272 6642 15328
rect 6698 15272 6703 15328
rect 4061 15270 6703 15272
rect 4061 15267 4127 15270
rect 6637 15267 6703 15270
rect 9121 15330 9187 15333
rect 11697 15330 11763 15333
rect 9121 15328 11763 15330
rect 9121 15272 9126 15328
rect 9182 15272 11702 15328
rect 11758 15272 11763 15328
rect 9121 15270 11763 15272
rect 9121 15267 9187 15270
rect 11697 15267 11763 15270
rect 3562 15264 3878 15265
rect 3562 15200 3568 15264
rect 3632 15200 3648 15264
rect 3712 15200 3728 15264
rect 3792 15200 3808 15264
rect 3872 15200 3878 15264
rect 3562 15199 3878 15200
rect 8562 15264 8878 15265
rect 8562 15200 8568 15264
rect 8632 15200 8648 15264
rect 8712 15200 8728 15264
rect 8792 15200 8808 15264
rect 8872 15200 8878 15264
rect 8562 15199 8878 15200
rect 6545 15194 6611 15197
rect 8385 15194 8451 15197
rect 6545 15192 8451 15194
rect 6545 15136 6550 15192
rect 6606 15136 8390 15192
rect 8446 15136 8451 15192
rect 6545 15134 8451 15136
rect 6545 15131 6611 15134
rect 8385 15131 8451 15134
rect 14000 15104 34000 15224
rect 16806 14959 16866 15104
rect 16757 14954 16866 14959
rect 105 14922 171 14925
rect 2773 14922 2839 14925
rect 105 14920 2839 14922
rect 105 14864 110 14920
rect 166 14864 2778 14920
rect 2834 14864 2839 14920
rect 105 14862 2839 14864
rect 105 14859 171 14862
rect 2773 14859 2839 14862
rect 8937 14922 9003 14925
rect 10685 14922 10751 14925
rect 8937 14920 10751 14922
rect 8937 14864 8942 14920
rect 8998 14864 10690 14920
rect 10746 14864 10751 14920
rect 16757 14898 16762 14954
rect 16818 14898 16866 14954
rect 16757 14896 16866 14898
rect 16757 14893 16823 14896
rect 8937 14862 10751 14864
rect 8937 14859 9003 14862
rect 10685 14859 10751 14862
rect 13813 14786 13879 14789
rect 14000 14786 34000 14816
rect 13813 14784 34000 14786
rect 13813 14728 13818 14784
rect 13874 14728 34000 14784
rect 13813 14726 34000 14728
rect 13813 14723 13879 14726
rect 2562 14720 2878 14721
rect 2562 14656 2568 14720
rect 2632 14656 2648 14720
rect 2712 14656 2728 14720
rect 2792 14656 2808 14720
rect 2872 14656 2878 14720
rect 2562 14655 2878 14656
rect 7562 14720 7878 14721
rect 7562 14656 7568 14720
rect 7632 14656 7648 14720
rect 7712 14656 7728 14720
rect 7792 14656 7808 14720
rect 7872 14656 7878 14720
rect 14000 14696 34000 14726
rect 7562 14655 7878 14656
rect 11053 14650 11119 14653
rect 11053 14648 13186 14650
rect 11053 14592 11058 14648
rect 11114 14592 13186 14648
rect 11053 14590 13186 14592
rect 11053 14587 11119 14590
rect 657 14514 723 14517
rect 4797 14514 4863 14517
rect 657 14512 4863 14514
rect 657 14456 662 14512
rect 718 14456 4802 14512
rect 4858 14456 4863 14512
rect 657 14454 4863 14456
rect 657 14451 723 14454
rect 4797 14451 4863 14454
rect 5441 14514 5507 14517
rect 12893 14514 12959 14517
rect 5441 14512 12959 14514
rect 5441 14456 5446 14512
rect 5502 14456 12898 14512
rect 12954 14456 12959 14512
rect 5441 14454 12959 14456
rect 5441 14451 5507 14454
rect 12893 14451 12959 14454
rect 565 14378 631 14381
rect 3601 14378 3667 14381
rect 565 14376 3667 14378
rect 565 14320 570 14376
rect 626 14320 3606 14376
rect 3662 14320 3667 14376
rect 565 14318 3667 14320
rect 565 14315 631 14318
rect 3601 14315 3667 14318
rect 7097 14378 7163 14381
rect 10317 14378 10383 14381
rect 7097 14376 10383 14378
rect 7097 14320 7102 14376
rect 7158 14320 10322 14376
rect 10378 14320 10383 14376
rect 7097 14318 10383 14320
rect 13126 14378 13186 14590
rect 14000 14378 34000 14408
rect 13126 14318 34000 14378
rect 7097 14315 7163 14318
rect 10317 14315 10383 14318
rect 14000 14288 34000 14318
rect 3562 14176 3878 14177
rect 3562 14112 3568 14176
rect 3632 14112 3648 14176
rect 3712 14112 3728 14176
rect 3792 14112 3808 14176
rect 3872 14112 3878 14176
rect 3562 14111 3878 14112
rect 8562 14176 8878 14177
rect 8562 14112 8568 14176
rect 8632 14112 8648 14176
rect 8712 14112 8728 14176
rect 8792 14112 8808 14176
rect 8872 14112 8878 14176
rect 8562 14111 8878 14112
rect 381 14106 447 14109
rect 2773 14106 2839 14109
rect 381 14104 2839 14106
rect 381 14048 386 14104
rect 442 14048 2778 14104
rect 2834 14048 2839 14104
rect 381 14046 2839 14048
rect 381 14043 447 14046
rect 2773 14043 2839 14046
rect 9305 14106 9371 14109
rect 11053 14106 11119 14109
rect 9305 14104 11119 14106
rect 9305 14048 9310 14104
rect 9366 14048 11058 14104
rect 11114 14048 11119 14104
rect 9305 14046 11119 14048
rect 9305 14043 9371 14046
rect 11053 14043 11119 14046
rect 2589 13970 2655 13973
rect 8017 13970 8083 13973
rect 2589 13968 8083 13970
rect 2589 13912 2594 13968
rect 2650 13912 8022 13968
rect 8078 13912 8083 13968
rect 2589 13910 8083 13912
rect 2589 13907 2655 13910
rect 8017 13907 8083 13910
rect 8937 13970 9003 13973
rect 13537 13970 13603 13973
rect 8937 13968 13603 13970
rect 8937 13912 8942 13968
rect 8998 13912 13542 13968
rect 13598 13912 13603 13968
rect 8937 13910 13603 13912
rect 8937 13907 9003 13910
rect 13537 13907 13603 13910
rect 13721 13970 13787 13973
rect 14000 13970 34000 14000
rect 13721 13968 34000 13970
rect 13721 13912 13726 13968
rect 13782 13912 34000 13968
rect 13721 13910 34000 13912
rect 13721 13907 13787 13910
rect 14000 13880 34000 13910
rect 289 13834 355 13837
rect 3049 13834 3115 13837
rect 289 13832 3115 13834
rect 289 13776 294 13832
rect 350 13776 3054 13832
rect 3110 13776 3115 13832
rect 289 13774 3115 13776
rect 289 13771 355 13774
rect 3049 13771 3115 13774
rect 4889 13834 4955 13837
rect 13445 13834 13511 13837
rect 4889 13832 13511 13834
rect 4889 13776 4894 13832
rect 4950 13776 13450 13832
rect 13506 13776 13511 13832
rect 4889 13774 13511 13776
rect 4889 13771 4955 13774
rect 13445 13771 13511 13774
rect 2562 13632 2878 13633
rect 2562 13568 2568 13632
rect 2632 13568 2648 13632
rect 2712 13568 2728 13632
rect 2792 13568 2808 13632
rect 2872 13568 2878 13632
rect 2562 13567 2878 13568
rect 7562 13632 7878 13633
rect 7562 13568 7568 13632
rect 7632 13568 7648 13632
rect 7712 13568 7728 13632
rect 7792 13568 7808 13632
rect 7872 13568 7878 13632
rect 7562 13567 7878 13568
rect 14000 13560 34000 13592
rect 14000 13504 15152 13560
rect 15208 13504 34000 13560
rect 14000 13472 34000 13504
rect 3509 13426 3575 13429
rect 5901 13426 5967 13429
rect 13629 13426 13695 13429
rect 3509 13424 5826 13426
rect 3509 13368 3514 13424
rect 3570 13368 5826 13424
rect 3509 13366 5826 13368
rect 3509 13363 3575 13366
rect 749 13290 815 13293
rect 4245 13290 4311 13293
rect 749 13288 4311 13290
rect 749 13232 754 13288
rect 810 13232 4250 13288
rect 4306 13232 4311 13288
rect 749 13230 4311 13232
rect 749 13227 815 13230
rect 4245 13227 4311 13230
rect 5766 13154 5826 13366
rect 5901 13424 13695 13426
rect 5901 13368 5906 13424
rect 5962 13368 13634 13424
rect 13690 13368 13695 13424
rect 5901 13366 13695 13368
rect 5901 13363 5967 13366
rect 13629 13363 13695 13366
rect 8109 13154 8175 13157
rect 5766 13152 8175 13154
rect 5766 13096 8114 13152
rect 8170 13096 8175 13152
rect 5766 13094 8175 13096
rect 8109 13091 8175 13094
rect 13813 13154 13879 13157
rect 14000 13154 34000 13184
rect 13813 13152 34000 13154
rect 13813 13096 13818 13152
rect 13874 13096 34000 13152
rect 13813 13094 34000 13096
rect 13813 13091 13879 13094
rect 3562 13088 3878 13089
rect 3562 13024 3568 13088
rect 3632 13024 3648 13088
rect 3712 13024 3728 13088
rect 3792 13024 3808 13088
rect 3872 13024 3878 13088
rect 3562 13023 3878 13024
rect 8562 13088 8878 13089
rect 8562 13024 8568 13088
rect 8632 13024 8648 13088
rect 8712 13024 8728 13088
rect 8792 13024 8808 13088
rect 8872 13024 8878 13088
rect 14000 13064 34000 13094
rect 8562 13023 8878 13024
rect 13 12882 79 12885
rect 3325 12882 3391 12885
rect 13 12880 3391 12882
rect 13 12824 18 12880
rect 74 12824 3330 12880
rect 3386 12824 3391 12880
rect 13 12822 3391 12824
rect 13 12819 79 12822
rect 3325 12819 3391 12822
rect 4337 12882 4403 12885
rect 7966 12882 7972 12884
rect 4337 12880 7972 12882
rect 4337 12824 4342 12880
rect 4398 12824 7972 12880
rect 4337 12822 7972 12824
rect 4337 12819 4403 12822
rect 7966 12820 7972 12822
rect 8036 12820 8042 12884
rect 8201 12882 8267 12885
rect 11789 12882 11855 12885
rect 8201 12880 11855 12882
rect 8201 12824 8206 12880
rect 8262 12824 11794 12880
rect 11850 12824 11855 12880
rect 8201 12822 11855 12824
rect 8201 12819 8267 12822
rect 11789 12819 11855 12822
rect 2589 12746 2655 12749
rect 11605 12746 11671 12749
rect 14000 12746 34000 12776
rect 2589 12744 11671 12746
rect 2589 12688 2594 12744
rect 2650 12688 11610 12744
rect 11666 12688 11671 12744
rect 2589 12686 11671 12688
rect 2589 12683 2655 12686
rect 11605 12683 11671 12686
rect 13862 12686 34000 12746
rect 3325 12610 3391 12613
rect 5533 12610 5599 12613
rect 3325 12608 5599 12610
rect 3325 12552 3330 12608
rect 3386 12552 5538 12608
rect 5594 12552 5599 12608
rect 3325 12550 5599 12552
rect 3325 12547 3391 12550
rect 5533 12547 5599 12550
rect 7966 12548 7972 12612
rect 8036 12610 8042 12612
rect 9305 12610 9371 12613
rect 8036 12608 9371 12610
rect 8036 12552 9310 12608
rect 9366 12552 9371 12608
rect 8036 12550 9371 12552
rect 8036 12548 8042 12550
rect 9305 12547 9371 12550
rect 11053 12610 11119 12613
rect 13169 12610 13235 12613
rect 11053 12608 13235 12610
rect 11053 12552 11058 12608
rect 11114 12552 13174 12608
rect 13230 12552 13235 12608
rect 11053 12550 13235 12552
rect 11053 12547 11119 12550
rect 13169 12547 13235 12550
rect 2562 12544 2878 12545
rect 2562 12480 2568 12544
rect 2632 12480 2648 12544
rect 2712 12480 2728 12544
rect 2792 12480 2808 12544
rect 2872 12480 2878 12544
rect 2562 12479 2878 12480
rect 7562 12544 7878 12545
rect 7562 12480 7568 12544
rect 7632 12480 7648 12544
rect 7712 12480 7728 12544
rect 7792 12480 7808 12544
rect 7872 12480 7878 12544
rect 7562 12479 7878 12480
rect 933 12476 999 12477
rect 933 12474 980 12476
rect 888 12472 980 12474
rect 888 12416 938 12472
rect 888 12414 980 12416
rect 933 12412 980 12414
rect 1044 12412 1050 12476
rect 1342 12412 1348 12476
rect 1412 12474 1418 12476
rect 1577 12474 1643 12477
rect 1412 12472 1643 12474
rect 1412 12416 1582 12472
rect 1638 12416 1643 12472
rect 1412 12414 1643 12416
rect 1412 12412 1418 12414
rect 933 12411 999 12412
rect 1577 12411 1643 12414
rect 13353 12474 13419 12477
rect 13862 12474 13922 12686
rect 14000 12656 34000 12686
rect 13353 12472 13922 12474
rect 13353 12416 13358 12472
rect 13414 12416 13922 12472
rect 13353 12414 13922 12416
rect 13353 12411 13419 12414
rect 4889 12338 4955 12341
rect 5993 12338 6059 12341
rect 8937 12338 9003 12341
rect 4889 12336 9003 12338
rect 4889 12280 4894 12336
rect 4950 12280 5998 12336
rect 6054 12280 8942 12336
rect 8998 12280 9003 12336
rect 4889 12278 9003 12280
rect 4889 12275 4955 12278
rect 5993 12275 6059 12278
rect 8937 12275 9003 12278
rect 14000 12336 34000 12368
rect 14000 12280 15152 12336
rect 15208 12280 34000 12336
rect 14000 12248 34000 12280
rect 5901 12202 5967 12205
rect 5901 12200 9138 12202
rect 5901 12144 5906 12200
rect 5962 12144 9138 12200
rect 5901 12142 9138 12144
rect 5901 12139 5967 12142
rect 4061 12066 4127 12069
rect 6913 12066 6979 12069
rect 4061 12064 6979 12066
rect 4061 12008 4066 12064
rect 4122 12008 6918 12064
rect 6974 12008 6979 12064
rect 4061 12006 6979 12008
rect 9078 12066 9138 12142
rect 12709 12066 12775 12069
rect 9078 12064 12775 12066
rect 9078 12008 12714 12064
rect 12770 12008 12775 12064
rect 9078 12006 12775 12008
rect 4061 12003 4127 12006
rect 6913 12003 6979 12006
rect 12709 12003 12775 12006
rect 3562 12000 3878 12001
rect 3562 11936 3568 12000
rect 3632 11936 3648 12000
rect 3712 11936 3728 12000
rect 3792 11936 3808 12000
rect 3872 11936 3878 12000
rect 3562 11935 3878 11936
rect 8562 12000 8878 12001
rect 8562 11936 8568 12000
rect 8632 11936 8648 12000
rect 8712 11936 8728 12000
rect 8792 11936 8808 12000
rect 8872 11936 8878 12000
rect 8562 11935 8878 11936
rect 11789 11930 11855 11933
rect 14000 11930 34000 11960
rect 11789 11928 34000 11930
rect 11789 11872 11794 11928
rect 11850 11872 34000 11928
rect 11789 11870 34000 11872
rect 11789 11867 11855 11870
rect 14000 11840 34000 11870
rect 8845 11794 8911 11797
rect 11881 11794 11947 11797
rect 8845 11792 11947 11794
rect 8845 11736 8850 11792
rect 8906 11736 11886 11792
rect 11942 11736 11947 11792
rect 8845 11734 11947 11736
rect 8845 11731 8911 11734
rect 11881 11731 11947 11734
rect 1485 11658 1551 11661
rect 4153 11658 4219 11661
rect 12801 11658 12867 11661
rect 1485 11656 4219 11658
rect 1485 11600 1490 11656
rect 1546 11600 4158 11656
rect 4214 11600 4219 11656
rect 1485 11598 4219 11600
rect 1485 11595 1551 11598
rect 4153 11595 4219 11598
rect 12390 11656 12867 11658
rect 12390 11600 12806 11656
rect 12862 11600 12867 11656
rect 12390 11598 12867 11600
rect 12390 11522 12450 11598
rect 12801 11595 12867 11598
rect 7974 11462 12450 11522
rect 14000 11520 34000 11552
rect 14000 11464 15152 11520
rect 15208 11464 34000 11520
rect 2562 11456 2878 11457
rect 2562 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2878 11456
rect 2562 11391 2878 11392
rect 7562 11456 7878 11457
rect 7562 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7878 11456
rect 7562 11391 7878 11392
rect 3417 11250 3483 11253
rect 7974 11250 8034 11462
rect 14000 11432 34000 11464
rect 8753 11386 8819 11389
rect 12525 11386 12591 11389
rect 8753 11384 12591 11386
rect 8753 11328 8758 11384
rect 8814 11328 12530 11384
rect 12586 11328 12591 11384
rect 8753 11326 12591 11328
rect 8753 11323 8819 11326
rect 12525 11323 12591 11326
rect 3417 11248 8034 11250
rect 3417 11192 3422 11248
rect 3478 11192 8034 11248
rect 3417 11190 8034 11192
rect 3417 11187 3483 11190
rect 197 11114 263 11117
rect 4153 11114 4219 11117
rect 197 11112 4219 11114
rect 197 11056 202 11112
rect 258 11056 4158 11112
rect 4214 11056 4219 11112
rect 197 11054 4219 11056
rect 197 11051 263 11054
rect 4153 11051 4219 11054
rect 4981 11114 5047 11117
rect 7005 11114 7071 11117
rect 4981 11112 7071 11114
rect 4981 11056 4986 11112
rect 5042 11056 7010 11112
rect 7066 11056 7071 11112
rect 4981 11054 7071 11056
rect 4981 11051 5047 11054
rect 7005 11051 7071 11054
rect 7189 11114 7255 11117
rect 13353 11114 13419 11117
rect 7189 11112 13419 11114
rect 7189 11056 7194 11112
rect 7250 11056 13358 11112
rect 13414 11056 13419 11112
rect 7189 11054 13419 11056
rect 7189 11051 7255 11054
rect 13353 11051 13419 11054
rect 13813 11114 13879 11117
rect 14000 11114 34000 11144
rect 13813 11112 34000 11114
rect 13813 11056 13818 11112
rect 13874 11056 34000 11112
rect 13813 11054 34000 11056
rect 13813 11051 13879 11054
rect 14000 11024 34000 11054
rect 3562 10912 3878 10913
rect 3562 10848 3568 10912
rect 3632 10848 3648 10912
rect 3712 10848 3728 10912
rect 3792 10848 3808 10912
rect 3872 10848 3878 10912
rect 3562 10847 3878 10848
rect 8562 10912 8878 10913
rect 8562 10848 8568 10912
rect 8632 10848 8648 10912
rect 8712 10848 8728 10912
rect 8792 10848 8808 10912
rect 8872 10848 8878 10912
rect 8562 10847 8878 10848
rect 9673 10842 9739 10845
rect 13813 10842 13879 10845
rect 9673 10840 13879 10842
rect 9673 10784 9678 10840
rect 9734 10784 13818 10840
rect 13874 10784 13879 10840
rect 9673 10782 13879 10784
rect 9673 10779 9739 10782
rect 13813 10779 13879 10782
rect 4889 10706 4955 10709
rect 9213 10706 9279 10709
rect 4889 10704 9279 10706
rect 4889 10648 4894 10704
rect 4950 10648 9218 10704
rect 9274 10648 9279 10704
rect 4889 10646 9279 10648
rect 4889 10643 4955 10646
rect 9213 10643 9279 10646
rect 13721 10706 13787 10709
rect 14000 10706 34000 10736
rect 13721 10704 34000 10706
rect 13721 10648 13726 10704
rect 13782 10648 34000 10704
rect 13721 10646 34000 10648
rect 13721 10643 13787 10646
rect 14000 10616 34000 10646
rect 2497 10570 2563 10573
rect 9489 10570 9555 10573
rect 2497 10568 9555 10570
rect 2497 10512 2502 10568
rect 2558 10512 9494 10568
rect 9550 10512 9555 10568
rect 2497 10510 9555 10512
rect 2497 10507 2563 10510
rect 9489 10507 9555 10510
rect 12433 10434 12499 10437
rect 12390 10432 12499 10434
rect 12390 10376 12438 10432
rect 12494 10376 12499 10432
rect 12390 10371 12499 10376
rect 2562 10368 2878 10369
rect 2562 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2878 10368
rect 2562 10303 2878 10304
rect 7562 10368 7878 10369
rect 7562 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7878 10368
rect 7562 10303 7878 10304
rect 3049 10298 3115 10301
rect 5717 10298 5783 10301
rect 3049 10296 5783 10298
rect 3049 10240 3054 10296
rect 3110 10240 5722 10296
rect 5778 10240 5783 10296
rect 3049 10238 5783 10240
rect 3049 10235 3115 10238
rect 5717 10235 5783 10238
rect 2037 10162 2103 10165
rect 5625 10162 5691 10165
rect 2037 10160 5691 10162
rect 2037 10104 2042 10160
rect 2098 10104 5630 10160
rect 5686 10104 5691 10160
rect 2037 10102 5691 10104
rect 2037 10099 2103 10102
rect 5625 10099 5691 10102
rect 5809 10162 5875 10165
rect 12390 10162 12450 10371
rect 14000 10296 34000 10328
rect 14000 10240 15152 10296
rect 15208 10240 34000 10296
rect 14000 10208 34000 10240
rect 5809 10160 12450 10162
rect 5809 10104 5814 10160
rect 5870 10104 12450 10160
rect 5809 10102 12450 10104
rect 5809 10099 5875 10102
rect 3141 10026 3207 10029
rect 4429 10026 4495 10029
rect 3141 10024 4495 10026
rect 3141 9968 3146 10024
rect 3202 9968 4434 10024
rect 4490 9968 4495 10024
rect 3141 9966 4495 9968
rect 3141 9963 3207 9966
rect 4429 9963 4495 9966
rect 8017 10026 8083 10029
rect 12617 10026 12683 10029
rect 8017 10024 12683 10026
rect 8017 9968 8022 10024
rect 8078 9968 12622 10024
rect 12678 9968 12683 10024
rect 8017 9966 12683 9968
rect 8017 9963 8083 9966
rect 12617 9963 12683 9966
rect 7005 9890 7071 9893
rect 8201 9890 8267 9893
rect 7005 9888 8267 9890
rect 7005 9832 7010 9888
rect 7066 9832 8206 9888
rect 8262 9832 8267 9888
rect 7005 9830 8267 9832
rect 7005 9827 7071 9830
rect 8201 9827 8267 9830
rect 9121 9890 9187 9893
rect 13077 9890 13143 9893
rect 9121 9888 13143 9890
rect 9121 9832 9126 9888
rect 9182 9832 13082 9888
rect 13138 9832 13143 9888
rect 9121 9830 13143 9832
rect 9121 9827 9187 9830
rect 13077 9827 13143 9830
rect 13813 9890 13879 9893
rect 14000 9890 34000 9920
rect 13813 9888 34000 9890
rect 13813 9832 13818 9888
rect 13874 9832 34000 9888
rect 13813 9830 34000 9832
rect 13813 9827 13879 9830
rect 3562 9824 3878 9825
rect 3562 9760 3568 9824
rect 3632 9760 3648 9824
rect 3712 9760 3728 9824
rect 3792 9760 3808 9824
rect 3872 9760 3878 9824
rect 3562 9759 3878 9760
rect 8562 9824 8878 9825
rect 8562 9760 8568 9824
rect 8632 9760 8648 9824
rect 8712 9760 8728 9824
rect 8792 9760 8808 9824
rect 8872 9760 8878 9824
rect 14000 9800 34000 9830
rect 8562 9759 8878 9760
rect 54 9692 60 9756
rect 124 9754 130 9756
rect 3233 9754 3299 9757
rect 124 9752 3299 9754
rect 124 9696 3238 9752
rect 3294 9696 3299 9752
rect 124 9694 3299 9696
rect 124 9692 130 9694
rect 3233 9691 3299 9694
rect 5993 9754 6059 9757
rect 8293 9754 8359 9757
rect 5993 9752 8359 9754
rect 5993 9696 5998 9752
rect 6054 9696 8298 9752
rect 8354 9696 8359 9752
rect 5993 9694 8359 9696
rect 5993 9691 6059 9694
rect 8293 9691 8359 9694
rect 5809 9618 5875 9621
rect 8937 9618 9003 9621
rect 5809 9616 9003 9618
rect 5809 9560 5814 9616
rect 5870 9560 8942 9616
rect 8998 9560 9003 9616
rect 5809 9558 9003 9560
rect 5809 9555 5875 9558
rect 8937 9555 9003 9558
rect 2681 9482 2747 9485
rect 11697 9482 11763 9485
rect 2681 9480 11763 9482
rect 2681 9424 2686 9480
rect 2742 9424 11702 9480
rect 11758 9424 11763 9480
rect 2681 9422 11763 9424
rect 2681 9419 2747 9422
rect 11697 9419 11763 9422
rect 13813 9482 13879 9485
rect 14000 9482 34000 9512
rect 13813 9480 34000 9482
rect 13813 9424 13818 9480
rect 13874 9424 34000 9480
rect 13813 9422 34000 9424
rect 13813 9419 13879 9422
rect 14000 9392 34000 9422
rect 4429 9346 4495 9349
rect 7005 9346 7071 9349
rect 4429 9344 7071 9346
rect 4429 9288 4434 9344
rect 4490 9288 7010 9344
rect 7066 9288 7071 9344
rect 4429 9286 7071 9288
rect 4429 9283 4495 9286
rect 7005 9283 7071 9286
rect 2562 9280 2878 9281
rect 2562 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2878 9280
rect 2562 9215 2878 9216
rect 7562 9280 7878 9281
rect 7562 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7878 9280
rect 7562 9215 7878 9216
rect 3049 9208 3115 9213
rect 3049 9152 3054 9208
rect 3110 9152 3115 9208
rect 3049 9147 3115 9152
rect 8017 9210 8083 9213
rect 10041 9210 10107 9213
rect 8017 9208 10107 9210
rect 8017 9152 8022 9208
rect 8078 9152 10046 9208
rect 10102 9152 10107 9208
rect 8017 9150 10107 9152
rect 8017 9147 8083 9150
rect 10041 9147 10107 9150
rect 3052 9074 3112 9147
rect 8334 9074 8340 9076
rect 3052 9014 8340 9074
rect 8334 9012 8340 9014
rect 8404 9012 8410 9076
rect 13813 9074 13879 9077
rect 14000 9074 34000 9104
rect 13813 9072 34000 9074
rect 13813 9016 13818 9072
rect 13874 9016 34000 9072
rect 13813 9014 34000 9016
rect 13813 9011 13879 9014
rect 14000 8984 34000 9014
rect 5349 8938 5415 8941
rect 8937 8938 9003 8941
rect 5349 8936 9003 8938
rect 5349 8880 5354 8936
rect 5410 8880 8942 8936
rect 8998 8880 9003 8936
rect 5349 8878 9003 8880
rect 5349 8875 5415 8878
rect 8937 8875 9003 8878
rect 5809 8802 5875 8805
rect 8017 8802 8083 8805
rect 5809 8800 8083 8802
rect 5809 8744 5814 8800
rect 5870 8744 8022 8800
rect 8078 8744 8083 8800
rect 5809 8742 8083 8744
rect 5809 8739 5875 8742
rect 8017 8739 8083 8742
rect 3562 8736 3878 8737
rect 3562 8672 3568 8736
rect 3632 8672 3648 8736
rect 3712 8672 3728 8736
rect 3792 8672 3808 8736
rect 3872 8672 3878 8736
rect 3562 8671 3878 8672
rect 8562 8736 8878 8737
rect 8562 8672 8568 8736
rect 8632 8672 8648 8736
rect 8712 8672 8728 8736
rect 8792 8672 8808 8736
rect 8872 8672 8878 8736
rect 8562 8671 8878 8672
rect 14000 8666 34000 8696
rect 9630 8606 34000 8666
rect 5625 8530 5691 8533
rect 9630 8530 9690 8606
rect 14000 8576 34000 8606
rect 5625 8528 9690 8530
rect 5625 8472 5630 8528
rect 5686 8472 9690 8528
rect 5625 8470 9690 8472
rect 5625 8467 5691 8470
rect 1117 8394 1183 8397
rect 2773 8394 2839 8397
rect 1117 8392 2839 8394
rect 1117 8336 1122 8392
rect 1178 8336 2778 8392
rect 2834 8336 2839 8392
rect 1117 8334 2839 8336
rect 1117 8331 1183 8334
rect 2773 8331 2839 8334
rect 3877 8394 3943 8397
rect 5901 8394 5967 8397
rect 3877 8392 5967 8394
rect 3877 8336 3882 8392
rect 3938 8336 5906 8392
rect 5962 8336 5967 8392
rect 3877 8334 5967 8336
rect 3877 8331 3943 8334
rect 5901 8331 5967 8334
rect 8201 8394 8267 8397
rect 12985 8394 13051 8397
rect 8201 8392 13051 8394
rect 8201 8336 8206 8392
rect 8262 8336 12990 8392
rect 13046 8336 13051 8392
rect 8201 8334 13051 8336
rect 8201 8331 8267 8334
rect 12985 8331 13051 8334
rect 3233 8258 3299 8261
rect 7097 8258 7163 8261
rect 3233 8256 7163 8258
rect 3233 8200 3238 8256
rect 3294 8200 7102 8256
rect 7158 8200 7163 8256
rect 3233 8198 7163 8200
rect 3233 8195 3299 8198
rect 7097 8195 7163 8198
rect 11789 8258 11855 8261
rect 14000 8258 34000 8288
rect 11789 8256 34000 8258
rect 11789 8200 11794 8256
rect 11850 8200 34000 8256
rect 11789 8198 34000 8200
rect 11789 8195 11855 8198
rect 2562 8192 2878 8193
rect 2562 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2878 8192
rect 2562 8127 2878 8128
rect 7562 8192 7878 8193
rect 7562 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7878 8192
rect 14000 8168 34000 8198
rect 7562 8127 7878 8128
rect 4102 8060 4108 8124
rect 4172 8122 4178 8124
rect 5165 8122 5231 8125
rect 4172 8120 5231 8122
rect 4172 8064 5170 8120
rect 5226 8064 5231 8120
rect 4172 8062 5231 8064
rect 4172 8060 4178 8062
rect 5165 8059 5231 8062
rect 2313 7850 2379 7853
rect 5533 7850 5599 7853
rect 2313 7848 5599 7850
rect 2313 7792 2318 7848
rect 2374 7792 5538 7848
rect 5594 7792 5599 7848
rect 2313 7790 5599 7792
rect 2313 7787 2379 7790
rect 5533 7787 5599 7790
rect 13721 7850 13787 7853
rect 14000 7850 34000 7880
rect 13721 7848 34000 7850
rect 13721 7792 13726 7848
rect 13782 7792 34000 7848
rect 13721 7790 34000 7792
rect 13721 7787 13787 7790
rect 14000 7760 34000 7790
rect 3562 7648 3878 7649
rect 3562 7584 3568 7648
rect 3632 7584 3648 7648
rect 3712 7584 3728 7648
rect 3792 7584 3808 7648
rect 3872 7584 3878 7648
rect 3562 7583 3878 7584
rect 8562 7648 8878 7649
rect 8562 7584 8568 7648
rect 8632 7584 8648 7648
rect 8712 7584 8728 7648
rect 8792 7584 8808 7648
rect 8872 7584 8878 7648
rect 8562 7583 8878 7584
rect 13261 7442 13327 7445
rect 14000 7442 34000 7472
rect 13261 7440 34000 7442
rect 13261 7384 13266 7440
rect 13322 7384 34000 7440
rect 13261 7382 34000 7384
rect 13261 7379 13327 7382
rect 14000 7352 34000 7382
rect 3233 7306 3299 7309
rect 3233 7304 8402 7306
rect 3233 7248 3238 7304
rect 3294 7248 8402 7304
rect 3233 7246 8402 7248
rect 3233 7243 3299 7246
rect 5533 7170 5599 7173
rect 7097 7170 7163 7173
rect 5533 7168 7163 7170
rect 5533 7112 5538 7168
rect 5594 7112 7102 7168
rect 7158 7112 7163 7168
rect 5533 7110 7163 7112
rect 5533 7107 5599 7110
rect 7097 7107 7163 7110
rect 2562 7104 2878 7105
rect 2562 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2878 7104
rect 2562 7039 2878 7040
rect 7562 7104 7878 7105
rect 7562 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7878 7104
rect 7562 7039 7878 7040
rect 4061 7034 4127 7037
rect 6361 7034 6427 7037
rect 4061 7032 6427 7034
rect 4061 6976 4066 7032
rect 4122 6976 6366 7032
rect 6422 6976 6427 7032
rect 4061 6974 6427 6976
rect 4061 6971 4127 6974
rect 6361 6971 6427 6974
rect 8342 6901 8402 7246
rect 11881 7034 11947 7037
rect 14000 7034 34000 7064
rect 11881 7032 34000 7034
rect 11881 6976 11886 7032
rect 11942 6976 34000 7032
rect 11881 6974 34000 6976
rect 11881 6971 11947 6974
rect 14000 6944 34000 6974
rect 5165 6898 5231 6901
rect 6269 6898 6335 6901
rect 5165 6896 6335 6898
rect 5165 6840 5170 6896
rect 5226 6840 6274 6896
rect 6330 6840 6335 6896
rect 5165 6838 6335 6840
rect 8342 6896 8451 6901
rect 8342 6840 8390 6896
rect 8446 6840 8451 6896
rect 8342 6838 8451 6840
rect 5165 6835 5231 6838
rect 6269 6835 6335 6838
rect 8385 6835 8451 6838
rect 5717 6762 5783 6765
rect 11789 6762 11855 6765
rect 5717 6760 11855 6762
rect 5717 6704 5722 6760
rect 5778 6704 11794 6760
rect 11850 6704 11855 6760
rect 5717 6702 11855 6704
rect 5717 6699 5783 6702
rect 11789 6699 11855 6702
rect 11237 6626 11303 6629
rect 14000 6626 34000 6656
rect 11237 6624 34000 6626
rect 11237 6568 11242 6624
rect 11298 6568 34000 6624
rect 11237 6566 34000 6568
rect 11237 6563 11303 6566
rect 3562 6560 3878 6561
rect 3562 6496 3568 6560
rect 3632 6496 3648 6560
rect 3712 6496 3728 6560
rect 3792 6496 3808 6560
rect 3872 6496 3878 6560
rect 3562 6495 3878 6496
rect 8562 6560 8878 6561
rect 8562 6496 8568 6560
rect 8632 6496 8648 6560
rect 8712 6496 8728 6560
rect 8792 6496 8808 6560
rect 8872 6496 8878 6560
rect 14000 6536 34000 6566
rect 8562 6495 8878 6496
rect 2405 6354 2471 6357
rect 13813 6354 13879 6357
rect 2405 6352 13879 6354
rect 2405 6296 2410 6352
rect 2466 6296 13818 6352
rect 13874 6296 13879 6352
rect 2405 6294 13879 6296
rect 2405 6291 2471 6294
rect 13813 6291 13879 6294
rect 6637 6218 6703 6221
rect 9121 6218 9187 6221
rect 6637 6216 9187 6218
rect 6637 6160 6642 6216
rect 6698 6160 9126 6216
rect 9182 6160 9187 6216
rect 6637 6158 9187 6160
rect 6637 6155 6703 6158
rect 9121 6155 9187 6158
rect 12341 6218 12407 6221
rect 12893 6218 12959 6221
rect 12341 6216 12959 6218
rect 12341 6160 12346 6216
rect 12402 6160 12898 6216
rect 12954 6160 12959 6216
rect 12341 6158 12959 6160
rect 12341 6155 12407 6158
rect 12893 6155 12959 6158
rect 13353 6218 13419 6221
rect 14000 6218 34000 6248
rect 13353 6216 34000 6218
rect 13353 6160 13358 6216
rect 13414 6160 34000 6216
rect 13353 6158 34000 6160
rect 13353 6155 13419 6158
rect 14000 6128 34000 6158
rect 3049 6082 3115 6085
rect 7189 6082 7255 6085
rect 3049 6080 7255 6082
rect 3049 6024 3054 6080
rect 3110 6024 7194 6080
rect 7250 6024 7255 6080
rect 3049 6022 7255 6024
rect 3049 6019 3115 6022
rect 7189 6019 7255 6022
rect 8201 6082 8267 6085
rect 10501 6082 10567 6085
rect 8201 6080 10567 6082
rect 8201 6024 8206 6080
rect 8262 6024 10506 6080
rect 10562 6024 10567 6080
rect 8201 6022 10567 6024
rect 8201 6019 8267 6022
rect 10501 6019 10567 6022
rect 2562 6016 2878 6017
rect 2562 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2878 6016
rect 2562 5951 2878 5952
rect 7562 6016 7878 6017
rect 7562 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7878 6016
rect 7562 5951 7878 5952
rect 5349 5946 5415 5949
rect 6177 5946 6243 5949
rect 5349 5944 6243 5946
rect 5349 5888 5354 5944
rect 5410 5888 6182 5944
rect 6238 5888 6243 5944
rect 5349 5886 6243 5888
rect 5349 5883 5415 5886
rect 6177 5883 6243 5886
rect 1945 5810 2011 5813
rect 4705 5810 4771 5813
rect 6545 5810 6611 5813
rect 1945 5808 6611 5810
rect 1945 5752 1950 5808
rect 2006 5752 4710 5808
rect 4766 5752 6550 5808
rect 6606 5752 6611 5808
rect 1945 5750 6611 5752
rect 1945 5747 2011 5750
rect 4705 5747 4771 5750
rect 6545 5747 6611 5750
rect 9673 5810 9739 5813
rect 13445 5810 13511 5813
rect 9673 5808 13511 5810
rect 9673 5752 9678 5808
rect 9734 5752 13450 5808
rect 13506 5752 13511 5808
rect 9673 5750 13511 5752
rect 9673 5747 9739 5750
rect 13445 5747 13511 5750
rect 13813 5810 13879 5813
rect 14000 5810 34000 5840
rect 13813 5808 34000 5810
rect 13813 5752 13818 5808
rect 13874 5752 34000 5808
rect 13813 5750 34000 5752
rect 13813 5747 13879 5750
rect 14000 5720 34000 5750
rect 13 5674 79 5677
rect 2497 5674 2563 5677
rect 13 5672 2563 5674
rect 13 5616 18 5672
rect 74 5616 2502 5672
rect 2558 5616 2563 5672
rect 13 5614 2563 5616
rect 13 5611 79 5614
rect 2497 5611 2563 5614
rect 3417 5674 3483 5677
rect 4337 5674 4403 5677
rect 3417 5672 4403 5674
rect 3417 5616 3422 5672
rect 3478 5616 4342 5672
rect 4398 5616 4403 5672
rect 3417 5614 4403 5616
rect 3417 5611 3483 5614
rect 4337 5611 4403 5614
rect 6177 5674 6243 5677
rect 8845 5674 8911 5677
rect 6177 5672 8911 5674
rect 6177 5616 6182 5672
rect 6238 5616 8850 5672
rect 8906 5616 8911 5672
rect 6177 5614 8911 5616
rect 6177 5611 6243 5614
rect 8845 5611 8911 5614
rect 11053 5674 11119 5677
rect 13537 5674 13603 5677
rect 11053 5672 13603 5674
rect 11053 5616 11058 5672
rect 11114 5616 13542 5672
rect 13598 5616 13603 5672
rect 11053 5614 13603 5616
rect 11053 5611 11119 5614
rect 13537 5611 13603 5614
rect 9857 5538 9923 5541
rect 12709 5538 12775 5541
rect 9857 5536 12775 5538
rect 9857 5480 9862 5536
rect 9918 5480 12714 5536
rect 12770 5480 12775 5536
rect 9857 5478 12775 5480
rect 9857 5475 9923 5478
rect 12709 5475 12775 5478
rect 3562 5472 3878 5473
rect 3562 5408 3568 5472
rect 3632 5408 3648 5472
rect 3712 5408 3728 5472
rect 3792 5408 3808 5472
rect 3872 5408 3878 5472
rect 3562 5407 3878 5408
rect 8562 5472 8878 5473
rect 8562 5408 8568 5472
rect 8632 5408 8648 5472
rect 8712 5408 8728 5472
rect 8792 5408 8808 5472
rect 8872 5408 8878 5472
rect 8562 5407 8878 5408
rect 2129 5402 2195 5405
rect 3325 5402 3391 5405
rect 2129 5400 3391 5402
rect 2129 5344 2134 5400
rect 2190 5344 3330 5400
rect 3386 5344 3391 5400
rect 2129 5342 3391 5344
rect 2129 5339 2195 5342
rect 3325 5339 3391 5342
rect 10317 5402 10383 5405
rect 14000 5402 34000 5432
rect 10317 5400 34000 5402
rect 10317 5344 10322 5400
rect 10378 5344 34000 5400
rect 10317 5342 34000 5344
rect 10317 5339 10383 5342
rect 14000 5312 34000 5342
rect 4889 5266 4955 5269
rect 11053 5266 11119 5269
rect 4889 5264 11119 5266
rect 4889 5208 4894 5264
rect 4950 5208 11058 5264
rect 11114 5208 11119 5264
rect 4889 5206 11119 5208
rect 4889 5203 4955 5206
rect 11053 5203 11119 5206
rect 11329 5266 11395 5269
rect 12525 5266 12591 5269
rect 11329 5264 12591 5266
rect 11329 5208 11334 5264
rect 11390 5208 12530 5264
rect 12586 5208 12591 5264
rect 11329 5206 12591 5208
rect 11329 5203 11395 5206
rect 12525 5203 12591 5206
rect 7189 5130 7255 5133
rect 9213 5130 9279 5133
rect 13721 5130 13787 5133
rect 7189 5128 8034 5130
rect 7189 5072 7194 5128
rect 7250 5072 8034 5128
rect 7189 5070 8034 5072
rect 7189 5067 7255 5070
rect 7562 4928 7878 4929
rect 7562 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7878 4928
rect 7562 4863 7878 4864
rect 5349 4858 5415 4861
rect 7281 4858 7347 4861
rect 5349 4856 7347 4858
rect 5349 4800 5354 4856
rect 5410 4800 7286 4856
rect 7342 4800 7347 4856
rect 5349 4798 7347 4800
rect 7974 4858 8034 5070
rect 9213 5128 13787 5130
rect 9213 5072 9218 5128
rect 9274 5072 13726 5128
rect 13782 5072 13787 5128
rect 9213 5070 13787 5072
rect 9213 5067 9279 5070
rect 13721 5067 13787 5070
rect 8569 4994 8635 4997
rect 12433 4994 12499 4997
rect 8569 4992 12499 4994
rect 8569 4936 8574 4992
rect 8630 4936 12438 4992
rect 12494 4936 12499 4992
rect 8569 4934 12499 4936
rect 8569 4931 8635 4934
rect 12433 4931 12499 4934
rect 12985 4994 13051 4997
rect 14000 4994 34000 5024
rect 12985 4992 34000 4994
rect 12985 4936 12990 4992
rect 13046 4936 34000 4992
rect 12985 4934 34000 4936
rect 12985 4931 13051 4934
rect 14000 4904 34000 4934
rect 13813 4858 13879 4861
rect 7974 4856 13879 4858
rect 7974 4800 13818 4856
rect 13874 4800 13879 4856
rect 7974 4798 13879 4800
rect 5349 4795 5415 4798
rect 7281 4795 7347 4798
rect 13813 4795 13879 4798
rect 1342 4660 1348 4724
rect 1412 4722 1418 4724
rect 3509 4722 3575 4725
rect 1412 4720 3575 4722
rect 1412 4664 3514 4720
rect 3570 4664 3575 4720
rect 1412 4662 3575 4664
rect 1412 4660 1418 4662
rect 3509 4659 3575 4662
rect 5993 4722 6059 4725
rect 11881 4722 11947 4725
rect 5993 4720 11947 4722
rect 5993 4664 5998 4720
rect 6054 4664 11886 4720
rect 11942 4664 11947 4720
rect 5993 4662 11947 4664
rect 5993 4659 6059 4662
rect 11881 4659 11947 4662
rect 1853 4586 1919 4589
rect 5717 4586 5783 4589
rect 1853 4584 5783 4586
rect 1853 4528 1858 4584
rect 1914 4528 5722 4584
rect 5778 4528 5783 4584
rect 1853 4526 5783 4528
rect 1853 4523 1919 4526
rect 5717 4523 5783 4526
rect 5993 4586 6059 4589
rect 9673 4586 9739 4589
rect 5993 4584 9739 4586
rect 5993 4528 5998 4584
rect 6054 4528 9678 4584
rect 9734 4528 9739 4584
rect 5993 4526 9739 4528
rect 5993 4523 6059 4526
rect 9673 4523 9739 4526
rect 11789 4586 11855 4589
rect 14000 4586 34000 4616
rect 11789 4584 34000 4586
rect 11789 4528 11794 4584
rect 11850 4528 34000 4584
rect 11789 4526 34000 4528
rect 11789 4523 11855 4526
rect 14000 4496 34000 4526
rect 4153 4450 4219 4453
rect 8201 4450 8267 4453
rect 4153 4448 8267 4450
rect 4153 4392 4158 4448
rect 4214 4392 8206 4448
rect 8262 4392 8267 4448
rect 4153 4390 8267 4392
rect 4153 4387 4219 4390
rect 8201 4387 8267 4390
rect 11053 4450 11119 4453
rect 13721 4450 13787 4453
rect 11053 4448 13787 4450
rect 11053 4392 11058 4448
rect 11114 4392 13726 4448
rect 13782 4392 13787 4448
rect 11053 4390 13787 4392
rect 11053 4387 11119 4390
rect 13721 4387 13787 4390
rect 3562 4384 3878 4385
rect 3562 4320 3568 4384
rect 3632 4320 3648 4384
rect 3712 4320 3728 4384
rect 3792 4320 3808 4384
rect 3872 4320 3878 4384
rect 3562 4319 3878 4320
rect 8562 4384 8878 4385
rect 8562 4320 8568 4384
rect 8632 4320 8648 4384
rect 8712 4320 8728 4384
rect 8792 4320 8808 4384
rect 8872 4320 8878 4384
rect 8562 4319 8878 4320
rect 14549 4314 14615 4317
rect 16297 4314 16363 4317
rect 14549 4312 16363 4314
rect 14549 4256 14554 4312
rect 14610 4256 16302 4312
rect 16358 4256 16363 4312
rect 14549 4254 16363 4256
rect 14549 4251 14615 4254
rect 16297 4251 16363 4254
rect 2405 4178 2471 4181
rect 4061 4178 4127 4181
rect 17033 4178 17099 4181
rect 2405 4176 2698 4178
rect 2405 4120 2410 4176
rect 2466 4120 2698 4176
rect 2405 4118 2698 4120
rect 2405 4115 2471 4118
rect 2638 4045 2698 4118
rect 4061 4176 17099 4178
rect 4061 4120 4066 4176
rect 4122 4120 17038 4176
rect 17094 4120 17099 4176
rect 4061 4118 17099 4120
rect 4061 4115 4127 4118
rect 17033 4115 17099 4118
rect 2405 4042 2471 4045
rect 2405 4040 2514 4042
rect 2405 3984 2410 4040
rect 2466 3984 2514 4040
rect 2405 3979 2514 3984
rect 2638 4040 2747 4045
rect 2638 3984 2686 4040
rect 2742 3984 2747 4040
rect 2638 3982 2747 3984
rect 2681 3979 2747 3982
rect 4061 4042 4127 4045
rect 16665 4042 16731 4045
rect 4061 4040 16731 4042
rect 4061 3984 4066 4040
rect 4122 3984 16670 4040
rect 16726 3984 16731 4040
rect 4061 3982 16731 3984
rect 4061 3979 4127 3982
rect 16665 3979 16731 3982
rect 2454 3400 2514 3979
rect 3325 3906 3391 3909
rect 6177 3906 6243 3909
rect 3325 3904 6243 3906
rect 3325 3848 3330 3904
rect 3386 3848 6182 3904
rect 6238 3848 6243 3904
rect 3325 3846 6243 3848
rect 3325 3843 3391 3846
rect 6177 3843 6243 3846
rect 9213 3906 9279 3909
rect 13261 3906 13327 3909
rect 9213 3904 13327 3906
rect 9213 3848 9218 3904
rect 9274 3848 13266 3904
rect 13322 3848 13327 3904
rect 9213 3846 13327 3848
rect 9213 3843 9279 3846
rect 13261 3843 13327 3846
rect 7562 3840 7878 3841
rect 7562 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7878 3840
rect 7562 3775 7878 3776
rect 2589 3770 2655 3773
rect 5441 3770 5507 3773
rect 2589 3768 5507 3770
rect 2589 3712 2594 3768
rect 2650 3712 5446 3768
rect 5502 3712 5507 3768
rect 2589 3710 5507 3712
rect 2589 3707 2655 3710
rect 5441 3707 5507 3710
rect 8201 3770 8267 3773
rect 12617 3770 12683 3773
rect 8201 3768 12683 3770
rect 8201 3712 8206 3768
rect 8262 3712 12622 3768
rect 12678 3712 12683 3768
rect 8201 3710 12683 3712
rect 8201 3707 8267 3710
rect 12617 3707 12683 3710
rect 2681 3634 2747 3637
rect 5625 3634 5691 3637
rect 2681 3632 5691 3634
rect 2681 3576 2686 3632
rect 2742 3576 5630 3632
rect 5686 3576 5691 3632
rect 2681 3574 5691 3576
rect 2681 3571 2747 3574
rect 5625 3571 5691 3574
rect 7005 3634 7071 3637
rect 11053 3634 11119 3637
rect 7005 3632 11119 3634
rect 7005 3576 7010 3632
rect 7066 3576 11058 3632
rect 11114 3576 11119 3632
rect 7005 3574 11119 3576
rect 7005 3571 7071 3574
rect 11053 3571 11119 3574
rect 11237 3634 11303 3637
rect 12801 3634 12867 3637
rect 11237 3632 12867 3634
rect 11237 3576 11242 3632
rect 11298 3576 12806 3632
rect 12862 3576 12867 3632
rect 11237 3574 12867 3576
rect 11237 3571 11303 3574
rect 12801 3571 12867 3574
rect 5993 3498 6059 3501
rect 10685 3498 10751 3501
rect 16113 3498 16179 3501
rect 5993 3496 9276 3498
rect 5993 3440 5998 3496
rect 6054 3440 9276 3496
rect 5993 3438 9276 3440
rect 5993 3435 6059 3438
rect 5073 3362 5139 3365
rect 8385 3362 8451 3365
rect 5073 3360 8451 3362
rect 5073 3304 5078 3360
rect 5134 3304 8390 3360
rect 8446 3304 8451 3360
rect 5073 3302 8451 3304
rect 9216 3362 9276 3438
rect 10685 3496 16179 3498
rect 10685 3440 10690 3496
rect 10746 3440 16118 3496
rect 16174 3440 16179 3496
rect 10685 3438 16179 3440
rect 10685 3435 10751 3438
rect 16113 3435 16179 3438
rect 13997 3362 14063 3365
rect 9216 3360 14063 3362
rect 9216 3304 14002 3360
rect 14058 3304 14063 3360
rect 9216 3302 14063 3304
rect 5073 3299 5139 3302
rect 8385 3299 8451 3302
rect 13997 3299 14063 3302
rect 3562 3296 3878 3297
rect 3562 3232 3568 3296
rect 3632 3232 3648 3296
rect 3712 3232 3728 3296
rect 3792 3232 3808 3296
rect 3872 3232 3878 3296
rect 3562 3231 3878 3232
rect 8562 3296 8878 3297
rect 8562 3232 8568 3296
rect 8632 3232 8648 3296
rect 8712 3232 8728 3296
rect 8792 3232 8808 3296
rect 8872 3232 8878 3296
rect 8562 3231 8878 3232
rect 9213 3226 9279 3229
rect 15837 3226 15903 3229
rect 9213 3224 15903 3226
rect 9213 3168 9218 3224
rect 9274 3168 15842 3224
rect 15898 3168 15903 3224
rect 9213 3166 15903 3168
rect 9213 3163 9279 3166
rect 15837 3163 15903 3166
rect 3141 3090 3207 3093
rect 4705 3090 4771 3093
rect 3141 3088 4771 3090
rect 3141 3032 3146 3088
rect 3202 3032 4710 3088
rect 4766 3032 4771 3088
rect 3141 3030 4771 3032
rect 3141 3027 3207 3030
rect 4705 3027 4771 3030
rect 5349 3090 5415 3093
rect 10869 3090 10935 3093
rect 5349 3088 10935 3090
rect 5349 3032 5354 3088
rect 5410 3032 10874 3088
rect 10930 3032 10935 3088
rect 5349 3030 10935 3032
rect 5349 3027 5415 3030
rect 10869 3027 10935 3030
rect 13169 2954 13235 2957
rect 7422 2952 13235 2954
rect 7422 2896 13174 2952
rect 13230 2896 13235 2952
rect 7422 2894 13235 2896
rect 4061 2684 4127 2685
rect 4061 2680 4108 2684
rect 4172 2682 4178 2684
rect 4061 2624 4066 2680
rect 4061 2620 4108 2624
rect 4172 2622 4218 2682
rect 4172 2620 4178 2622
rect 4061 2619 4127 2620
rect 2405 2546 2471 2549
rect 5625 2546 5691 2549
rect 2405 2544 5691 2546
rect 2405 2488 2410 2544
rect 2466 2488 5630 2544
rect 5686 2488 5691 2544
rect 2405 2486 5691 2488
rect 2405 2483 2471 2486
rect 5625 2483 5691 2486
rect 6085 2546 6151 2549
rect 7422 2546 7482 2894
rect 13169 2891 13235 2894
rect 8017 2818 8083 2821
rect 14549 2818 14615 2821
rect 8017 2816 14615 2818
rect 8017 2760 8022 2816
rect 8078 2760 14554 2816
rect 14610 2760 14615 2816
rect 8017 2758 14615 2760
rect 8017 2755 8083 2758
rect 14549 2755 14615 2758
rect 7562 2752 7878 2753
rect 7562 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7878 2752
rect 7562 2687 7878 2688
rect 8017 2682 8083 2685
rect 16573 2682 16639 2685
rect 8017 2680 16639 2682
rect 8017 2624 8022 2680
rect 8078 2624 16578 2680
rect 16634 2624 16639 2680
rect 8017 2622 16639 2624
rect 8017 2619 8083 2622
rect 16573 2619 16639 2622
rect 6085 2544 7482 2546
rect 6085 2488 6090 2544
rect 6146 2488 7482 2544
rect 6085 2486 7482 2488
rect 6085 2483 6151 2486
rect 8334 2484 8340 2548
rect 8404 2546 8410 2548
rect 8477 2546 8543 2549
rect 8404 2544 8543 2546
rect 8404 2488 8482 2544
rect 8538 2488 8543 2544
rect 8404 2486 8543 2488
rect 8404 2484 8410 2486
rect 8477 2483 8543 2486
rect 5625 2410 5691 2413
rect 10685 2410 10751 2413
rect 5625 2408 10751 2410
rect 5625 2352 5630 2408
rect 5686 2352 10690 2408
rect 10746 2352 10751 2408
rect 5625 2350 10751 2352
rect 5625 2347 5691 2350
rect 10685 2347 10751 2350
rect 3562 2208 3878 2209
rect 3562 2144 3568 2208
rect 3632 2144 3648 2208
rect 3712 2144 3728 2208
rect 3792 2144 3808 2208
rect 3872 2144 3878 2208
rect 3562 2143 3878 2144
rect 8562 2208 8878 2209
rect 8562 2144 8568 2208
rect 8632 2144 8648 2208
rect 8712 2144 8728 2208
rect 8792 2144 8808 2208
rect 8872 2144 8878 2208
rect 8562 2143 8878 2144
rect 6269 2002 6335 2005
rect 15285 2002 15351 2005
rect 6269 2000 15351 2002
rect 6269 1944 6274 2000
rect 6330 1944 15290 2000
rect 15346 1944 15351 2000
rect 6269 1942 15351 1944
rect 6269 1939 6335 1942
rect 15285 1939 15351 1942
rect 8477 1866 8543 1869
rect 11789 1866 11855 1869
rect 8477 1864 11855 1866
rect 8477 1808 8482 1864
rect 8538 1808 11794 1864
rect 11850 1808 11855 1864
rect 8477 1806 11855 1808
rect 8477 1803 8543 1806
rect 11789 1803 11855 1806
rect 2405 1730 2471 1733
rect 6545 1730 6611 1733
rect 2405 1728 6611 1730
rect 2405 1672 2410 1728
rect 2466 1672 6550 1728
rect 6606 1672 6611 1728
rect 2405 1670 6611 1672
rect 2405 1667 2471 1670
rect 6545 1667 6611 1670
rect 8661 1730 8727 1733
rect 10317 1730 10383 1733
rect 8661 1728 10383 1730
rect 8661 1672 8666 1728
rect 8722 1672 10322 1728
rect 10378 1672 10383 1728
rect 8661 1670 10383 1672
rect 8661 1667 8727 1670
rect 10317 1667 10383 1670
rect 7562 1664 7878 1665
rect 7562 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7878 1664
rect 7562 1599 7878 1600
rect 105 1596 171 1597
rect 54 1594 60 1596
rect 14 1534 60 1594
rect 124 1592 171 1596
rect 166 1536 171 1592
rect 54 1532 60 1534
rect 124 1532 171 1536
rect 105 1531 171 1532
rect 473 1594 539 1597
rect 1853 1594 1919 1597
rect 473 1592 1919 1594
rect 473 1536 478 1592
rect 534 1536 1858 1592
rect 1914 1536 1919 1592
rect 473 1534 1919 1536
rect 473 1531 539 1534
rect 1853 1531 1919 1534
rect 2313 1594 2379 1597
rect 4153 1594 4219 1597
rect 2313 1592 4219 1594
rect 2313 1536 2318 1592
rect 2374 1536 4158 1592
rect 4214 1536 4219 1592
rect 2313 1534 4219 1536
rect 2313 1531 2379 1534
rect 4153 1531 4219 1534
rect 5441 1594 5507 1597
rect 5441 1592 7482 1594
rect 5441 1536 5446 1592
rect 5502 1536 7482 1592
rect 5441 1534 7482 1536
rect 5441 1531 5507 1534
rect 197 1458 263 1461
rect 2773 1458 2839 1461
rect 197 1456 2839 1458
rect 197 1400 202 1456
rect 258 1400 2778 1456
rect 2834 1400 2839 1456
rect 197 1398 2839 1400
rect 197 1395 263 1398
rect 2773 1395 2839 1398
rect 2957 1458 3023 1461
rect 6821 1458 6887 1461
rect 2957 1456 6887 1458
rect 2957 1400 2962 1456
rect 3018 1400 6826 1456
rect 6882 1400 6887 1456
rect 2957 1398 6887 1400
rect 7422 1458 7482 1534
rect 12341 1458 12407 1461
rect 7422 1456 12407 1458
rect 7422 1400 12346 1456
rect 12402 1400 12407 1456
rect 7422 1398 12407 1400
rect 2957 1395 3023 1398
rect 6821 1395 6887 1398
rect 12341 1395 12407 1398
rect 1117 1322 1183 1325
rect 3601 1322 3667 1325
rect 1117 1320 3667 1322
rect 1117 1264 1122 1320
rect 1178 1264 3606 1320
rect 3662 1264 3667 1320
rect 1117 1262 3667 1264
rect 1117 1259 1183 1262
rect 3601 1259 3667 1262
rect 4061 1322 4127 1325
rect 7373 1322 7439 1325
rect 10777 1322 10843 1325
rect 4061 1320 7439 1322
rect 4061 1264 4066 1320
rect 4122 1264 7378 1320
rect 7434 1264 7439 1320
rect 4061 1262 7439 1264
rect 4061 1259 4127 1262
rect 7373 1259 7439 1262
rect 8342 1320 10843 1322
rect 8342 1264 10782 1320
rect 10838 1264 10843 1320
rect 8342 1262 10843 1264
rect 565 1186 631 1189
rect 3417 1186 3483 1189
rect 565 1184 3483 1186
rect 565 1128 570 1184
rect 626 1128 3422 1184
rect 3478 1128 3483 1184
rect 565 1126 3483 1128
rect 565 1123 631 1126
rect 3417 1123 3483 1126
rect 3562 1120 3878 1121
rect 3562 1056 3568 1120
rect 3632 1056 3648 1120
rect 3712 1056 3728 1120
rect 3792 1056 3808 1120
rect 3872 1056 3878 1120
rect 3562 1055 3878 1056
rect 381 914 447 917
rect 4705 914 4771 917
rect 381 912 4771 914
rect 381 856 386 912
rect 442 856 4710 912
rect 4766 856 4771 912
rect 381 854 4771 856
rect 381 851 447 854
rect 4705 851 4771 854
rect 4889 914 4955 917
rect 8342 914 8402 1262
rect 10777 1259 10843 1262
rect 8562 1120 8878 1121
rect 8562 1056 8568 1120
rect 8632 1056 8648 1120
rect 8712 1056 8728 1120
rect 8792 1056 8808 1120
rect 8872 1056 8878 1120
rect 8562 1055 8878 1056
rect 4889 912 8402 914
rect 4889 856 4894 912
rect 4950 856 8402 912
rect 4889 854 8402 856
rect 11697 914 11763 917
rect 16389 914 16455 917
rect 11697 912 16455 914
rect 11697 856 11702 912
rect 11758 856 16394 912
rect 16450 856 16455 912
rect 11697 854 16455 856
rect 4889 851 4955 854
rect 11697 851 11763 854
rect 16389 851 16455 854
rect 4337 778 4403 781
rect 7097 778 7163 781
rect 4337 776 7163 778
rect 4337 720 4342 776
rect 4398 720 7102 776
rect 7158 720 7163 776
rect 4337 718 7163 720
rect 4337 715 4403 718
rect 7097 715 7163 718
rect 7281 778 7347 781
rect 16481 778 16547 781
rect 7281 776 16547 778
rect 7281 720 7286 776
rect 7342 720 16486 776
rect 16542 720 16547 776
rect 7281 718 16547 720
rect 7281 715 7347 718
rect 16481 715 16547 718
rect 6729 642 6795 645
rect 16849 642 16915 645
rect 6729 640 16915 642
rect 6729 584 6734 640
rect 6790 584 16854 640
rect 16910 584 16915 640
rect 6729 582 16915 584
rect 6729 579 6795 582
rect 16849 579 16915 582
rect 6637 506 6703 509
rect 6913 506 6979 509
rect 6637 504 6979 506
rect 6637 448 6642 504
rect 6698 448 6918 504
rect 6974 448 6979 504
rect 6637 446 6979 448
rect 6637 443 6703 446
rect 6913 443 6979 446
rect 7097 506 7163 509
rect 11697 506 11763 509
rect 7097 504 11763 506
rect 7097 448 7102 504
rect 7158 448 11702 504
rect 11758 448 11763 504
rect 7097 446 11763 448
rect 7097 443 7163 446
rect 11697 443 11763 446
rect 4153 370 4219 373
rect 16757 370 16823 373
rect 4153 368 16823 370
rect 4153 312 4158 368
rect 4214 312 16762 368
rect 16818 312 16823 368
rect 4153 310 16823 312
rect 4153 307 4219 310
rect 16757 307 16823 310
rect 6913 234 6979 237
rect 11145 234 11211 237
rect 6913 232 11211 234
rect 6913 176 6918 232
rect 6974 176 11150 232
rect 11206 176 11211 232
rect 6913 174 11211 176
rect 6913 171 6979 174
rect 11145 171 11211 174
<< via3 >>
rect 2568 15804 2632 15808
rect 2568 15748 2572 15804
rect 2572 15748 2628 15804
rect 2628 15748 2632 15804
rect 2568 15744 2632 15748
rect 2648 15804 2712 15808
rect 2648 15748 2652 15804
rect 2652 15748 2708 15804
rect 2708 15748 2712 15804
rect 2648 15744 2712 15748
rect 2728 15804 2792 15808
rect 2728 15748 2732 15804
rect 2732 15748 2788 15804
rect 2788 15748 2792 15804
rect 2728 15744 2792 15748
rect 2808 15804 2872 15808
rect 2808 15748 2812 15804
rect 2812 15748 2868 15804
rect 2868 15748 2872 15804
rect 2808 15744 2872 15748
rect 7568 15804 7632 15808
rect 7568 15748 7572 15804
rect 7572 15748 7628 15804
rect 7628 15748 7632 15804
rect 7568 15744 7632 15748
rect 7648 15804 7712 15808
rect 7648 15748 7652 15804
rect 7652 15748 7708 15804
rect 7708 15748 7712 15804
rect 7648 15744 7712 15748
rect 7728 15804 7792 15808
rect 7728 15748 7732 15804
rect 7732 15748 7788 15804
rect 7788 15748 7792 15804
rect 7728 15744 7792 15748
rect 7808 15804 7872 15808
rect 7808 15748 7812 15804
rect 7812 15748 7868 15804
rect 7868 15748 7872 15804
rect 7808 15744 7872 15748
rect 980 15268 1044 15332
rect 3568 15260 3632 15264
rect 3568 15204 3572 15260
rect 3572 15204 3628 15260
rect 3628 15204 3632 15260
rect 3568 15200 3632 15204
rect 3648 15260 3712 15264
rect 3648 15204 3652 15260
rect 3652 15204 3708 15260
rect 3708 15204 3712 15260
rect 3648 15200 3712 15204
rect 3728 15260 3792 15264
rect 3728 15204 3732 15260
rect 3732 15204 3788 15260
rect 3788 15204 3792 15260
rect 3728 15200 3792 15204
rect 3808 15260 3872 15264
rect 3808 15204 3812 15260
rect 3812 15204 3868 15260
rect 3868 15204 3872 15260
rect 3808 15200 3872 15204
rect 8568 15260 8632 15264
rect 8568 15204 8572 15260
rect 8572 15204 8628 15260
rect 8628 15204 8632 15260
rect 8568 15200 8632 15204
rect 8648 15260 8712 15264
rect 8648 15204 8652 15260
rect 8652 15204 8708 15260
rect 8708 15204 8712 15260
rect 8648 15200 8712 15204
rect 8728 15260 8792 15264
rect 8728 15204 8732 15260
rect 8732 15204 8788 15260
rect 8788 15204 8792 15260
rect 8728 15200 8792 15204
rect 8808 15260 8872 15264
rect 8808 15204 8812 15260
rect 8812 15204 8868 15260
rect 8868 15204 8872 15260
rect 8808 15200 8872 15204
rect 2568 14716 2632 14720
rect 2568 14660 2572 14716
rect 2572 14660 2628 14716
rect 2628 14660 2632 14716
rect 2568 14656 2632 14660
rect 2648 14716 2712 14720
rect 2648 14660 2652 14716
rect 2652 14660 2708 14716
rect 2708 14660 2712 14716
rect 2648 14656 2712 14660
rect 2728 14716 2792 14720
rect 2728 14660 2732 14716
rect 2732 14660 2788 14716
rect 2788 14660 2792 14716
rect 2728 14656 2792 14660
rect 2808 14716 2872 14720
rect 2808 14660 2812 14716
rect 2812 14660 2868 14716
rect 2868 14660 2872 14716
rect 2808 14656 2872 14660
rect 7568 14716 7632 14720
rect 7568 14660 7572 14716
rect 7572 14660 7628 14716
rect 7628 14660 7632 14716
rect 7568 14656 7632 14660
rect 7648 14716 7712 14720
rect 7648 14660 7652 14716
rect 7652 14660 7708 14716
rect 7708 14660 7712 14716
rect 7648 14656 7712 14660
rect 7728 14716 7792 14720
rect 7728 14660 7732 14716
rect 7732 14660 7788 14716
rect 7788 14660 7792 14716
rect 7728 14656 7792 14660
rect 7808 14716 7872 14720
rect 7808 14660 7812 14716
rect 7812 14660 7868 14716
rect 7868 14660 7872 14716
rect 7808 14656 7872 14660
rect 3568 14172 3632 14176
rect 3568 14116 3572 14172
rect 3572 14116 3628 14172
rect 3628 14116 3632 14172
rect 3568 14112 3632 14116
rect 3648 14172 3712 14176
rect 3648 14116 3652 14172
rect 3652 14116 3708 14172
rect 3708 14116 3712 14172
rect 3648 14112 3712 14116
rect 3728 14172 3792 14176
rect 3728 14116 3732 14172
rect 3732 14116 3788 14172
rect 3788 14116 3792 14172
rect 3728 14112 3792 14116
rect 3808 14172 3872 14176
rect 3808 14116 3812 14172
rect 3812 14116 3868 14172
rect 3868 14116 3872 14172
rect 3808 14112 3872 14116
rect 8568 14172 8632 14176
rect 8568 14116 8572 14172
rect 8572 14116 8628 14172
rect 8628 14116 8632 14172
rect 8568 14112 8632 14116
rect 8648 14172 8712 14176
rect 8648 14116 8652 14172
rect 8652 14116 8708 14172
rect 8708 14116 8712 14172
rect 8648 14112 8712 14116
rect 8728 14172 8792 14176
rect 8728 14116 8732 14172
rect 8732 14116 8788 14172
rect 8788 14116 8792 14172
rect 8728 14112 8792 14116
rect 8808 14172 8872 14176
rect 8808 14116 8812 14172
rect 8812 14116 8868 14172
rect 8868 14116 8872 14172
rect 8808 14112 8872 14116
rect 2568 13628 2632 13632
rect 2568 13572 2572 13628
rect 2572 13572 2628 13628
rect 2628 13572 2632 13628
rect 2568 13568 2632 13572
rect 2648 13628 2712 13632
rect 2648 13572 2652 13628
rect 2652 13572 2708 13628
rect 2708 13572 2712 13628
rect 2648 13568 2712 13572
rect 2728 13628 2792 13632
rect 2728 13572 2732 13628
rect 2732 13572 2788 13628
rect 2788 13572 2792 13628
rect 2728 13568 2792 13572
rect 2808 13628 2872 13632
rect 2808 13572 2812 13628
rect 2812 13572 2868 13628
rect 2868 13572 2872 13628
rect 2808 13568 2872 13572
rect 7568 13628 7632 13632
rect 7568 13572 7572 13628
rect 7572 13572 7628 13628
rect 7628 13572 7632 13628
rect 7568 13568 7632 13572
rect 7648 13628 7712 13632
rect 7648 13572 7652 13628
rect 7652 13572 7708 13628
rect 7708 13572 7712 13628
rect 7648 13568 7712 13572
rect 7728 13628 7792 13632
rect 7728 13572 7732 13628
rect 7732 13572 7788 13628
rect 7788 13572 7792 13628
rect 7728 13568 7792 13572
rect 7808 13628 7872 13632
rect 7808 13572 7812 13628
rect 7812 13572 7868 13628
rect 7868 13572 7872 13628
rect 7808 13568 7872 13572
rect 3568 13084 3632 13088
rect 3568 13028 3572 13084
rect 3572 13028 3628 13084
rect 3628 13028 3632 13084
rect 3568 13024 3632 13028
rect 3648 13084 3712 13088
rect 3648 13028 3652 13084
rect 3652 13028 3708 13084
rect 3708 13028 3712 13084
rect 3648 13024 3712 13028
rect 3728 13084 3792 13088
rect 3728 13028 3732 13084
rect 3732 13028 3788 13084
rect 3788 13028 3792 13084
rect 3728 13024 3792 13028
rect 3808 13084 3872 13088
rect 3808 13028 3812 13084
rect 3812 13028 3868 13084
rect 3868 13028 3872 13084
rect 3808 13024 3872 13028
rect 8568 13084 8632 13088
rect 8568 13028 8572 13084
rect 8572 13028 8628 13084
rect 8628 13028 8632 13084
rect 8568 13024 8632 13028
rect 8648 13084 8712 13088
rect 8648 13028 8652 13084
rect 8652 13028 8708 13084
rect 8708 13028 8712 13084
rect 8648 13024 8712 13028
rect 8728 13084 8792 13088
rect 8728 13028 8732 13084
rect 8732 13028 8788 13084
rect 8788 13028 8792 13084
rect 8728 13024 8792 13028
rect 8808 13084 8872 13088
rect 8808 13028 8812 13084
rect 8812 13028 8868 13084
rect 8868 13028 8872 13084
rect 8808 13024 8872 13028
rect 7972 12820 8036 12884
rect 7972 12548 8036 12612
rect 2568 12540 2632 12544
rect 2568 12484 2572 12540
rect 2572 12484 2628 12540
rect 2628 12484 2632 12540
rect 2568 12480 2632 12484
rect 2648 12540 2712 12544
rect 2648 12484 2652 12540
rect 2652 12484 2708 12540
rect 2708 12484 2712 12540
rect 2648 12480 2712 12484
rect 2728 12540 2792 12544
rect 2728 12484 2732 12540
rect 2732 12484 2788 12540
rect 2788 12484 2792 12540
rect 2728 12480 2792 12484
rect 2808 12540 2872 12544
rect 2808 12484 2812 12540
rect 2812 12484 2868 12540
rect 2868 12484 2872 12540
rect 2808 12480 2872 12484
rect 7568 12540 7632 12544
rect 7568 12484 7572 12540
rect 7572 12484 7628 12540
rect 7628 12484 7632 12540
rect 7568 12480 7632 12484
rect 7648 12540 7712 12544
rect 7648 12484 7652 12540
rect 7652 12484 7708 12540
rect 7708 12484 7712 12540
rect 7648 12480 7712 12484
rect 7728 12540 7792 12544
rect 7728 12484 7732 12540
rect 7732 12484 7788 12540
rect 7788 12484 7792 12540
rect 7728 12480 7792 12484
rect 7808 12540 7872 12544
rect 7808 12484 7812 12540
rect 7812 12484 7868 12540
rect 7868 12484 7872 12540
rect 7808 12480 7872 12484
rect 980 12472 1044 12476
rect 980 12416 994 12472
rect 994 12416 1044 12472
rect 980 12412 1044 12416
rect 1348 12412 1412 12476
rect 3568 11996 3632 12000
rect 3568 11940 3572 11996
rect 3572 11940 3628 11996
rect 3628 11940 3632 11996
rect 3568 11936 3632 11940
rect 3648 11996 3712 12000
rect 3648 11940 3652 11996
rect 3652 11940 3708 11996
rect 3708 11940 3712 11996
rect 3648 11936 3712 11940
rect 3728 11996 3792 12000
rect 3728 11940 3732 11996
rect 3732 11940 3788 11996
rect 3788 11940 3792 11996
rect 3728 11936 3792 11940
rect 3808 11996 3872 12000
rect 3808 11940 3812 11996
rect 3812 11940 3868 11996
rect 3868 11940 3872 11996
rect 3808 11936 3872 11940
rect 8568 11996 8632 12000
rect 8568 11940 8572 11996
rect 8572 11940 8628 11996
rect 8628 11940 8632 11996
rect 8568 11936 8632 11940
rect 8648 11996 8712 12000
rect 8648 11940 8652 11996
rect 8652 11940 8708 11996
rect 8708 11940 8712 11996
rect 8648 11936 8712 11940
rect 8728 11996 8792 12000
rect 8728 11940 8732 11996
rect 8732 11940 8788 11996
rect 8788 11940 8792 11996
rect 8728 11936 8792 11940
rect 8808 11996 8872 12000
rect 8808 11940 8812 11996
rect 8812 11940 8868 11996
rect 8868 11940 8872 11996
rect 8808 11936 8872 11940
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 7568 11452 7632 11456
rect 7568 11396 7572 11452
rect 7572 11396 7628 11452
rect 7628 11396 7632 11452
rect 7568 11392 7632 11396
rect 7648 11452 7712 11456
rect 7648 11396 7652 11452
rect 7652 11396 7708 11452
rect 7708 11396 7712 11452
rect 7648 11392 7712 11396
rect 7728 11452 7792 11456
rect 7728 11396 7732 11452
rect 7732 11396 7788 11452
rect 7788 11396 7792 11452
rect 7728 11392 7792 11396
rect 7808 11452 7872 11456
rect 7808 11396 7812 11452
rect 7812 11396 7868 11452
rect 7868 11396 7872 11452
rect 7808 11392 7872 11396
rect 3568 10908 3632 10912
rect 3568 10852 3572 10908
rect 3572 10852 3628 10908
rect 3628 10852 3632 10908
rect 3568 10848 3632 10852
rect 3648 10908 3712 10912
rect 3648 10852 3652 10908
rect 3652 10852 3708 10908
rect 3708 10852 3712 10908
rect 3648 10848 3712 10852
rect 3728 10908 3792 10912
rect 3728 10852 3732 10908
rect 3732 10852 3788 10908
rect 3788 10852 3792 10908
rect 3728 10848 3792 10852
rect 3808 10908 3872 10912
rect 3808 10852 3812 10908
rect 3812 10852 3868 10908
rect 3868 10852 3872 10908
rect 3808 10848 3872 10852
rect 8568 10908 8632 10912
rect 8568 10852 8572 10908
rect 8572 10852 8628 10908
rect 8628 10852 8632 10908
rect 8568 10848 8632 10852
rect 8648 10908 8712 10912
rect 8648 10852 8652 10908
rect 8652 10852 8708 10908
rect 8708 10852 8712 10908
rect 8648 10848 8712 10852
rect 8728 10908 8792 10912
rect 8728 10852 8732 10908
rect 8732 10852 8788 10908
rect 8788 10852 8792 10908
rect 8728 10848 8792 10852
rect 8808 10908 8872 10912
rect 8808 10852 8812 10908
rect 8812 10852 8868 10908
rect 8868 10852 8872 10908
rect 8808 10848 8872 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 7568 10364 7632 10368
rect 7568 10308 7572 10364
rect 7572 10308 7628 10364
rect 7628 10308 7632 10364
rect 7568 10304 7632 10308
rect 7648 10364 7712 10368
rect 7648 10308 7652 10364
rect 7652 10308 7708 10364
rect 7708 10308 7712 10364
rect 7648 10304 7712 10308
rect 7728 10364 7792 10368
rect 7728 10308 7732 10364
rect 7732 10308 7788 10364
rect 7788 10308 7792 10364
rect 7728 10304 7792 10308
rect 7808 10364 7872 10368
rect 7808 10308 7812 10364
rect 7812 10308 7868 10364
rect 7868 10308 7872 10364
rect 7808 10304 7872 10308
rect 3568 9820 3632 9824
rect 3568 9764 3572 9820
rect 3572 9764 3628 9820
rect 3628 9764 3632 9820
rect 3568 9760 3632 9764
rect 3648 9820 3712 9824
rect 3648 9764 3652 9820
rect 3652 9764 3708 9820
rect 3708 9764 3712 9820
rect 3648 9760 3712 9764
rect 3728 9820 3792 9824
rect 3728 9764 3732 9820
rect 3732 9764 3788 9820
rect 3788 9764 3792 9820
rect 3728 9760 3792 9764
rect 3808 9820 3872 9824
rect 3808 9764 3812 9820
rect 3812 9764 3868 9820
rect 3868 9764 3872 9820
rect 3808 9760 3872 9764
rect 8568 9820 8632 9824
rect 8568 9764 8572 9820
rect 8572 9764 8628 9820
rect 8628 9764 8632 9820
rect 8568 9760 8632 9764
rect 8648 9820 8712 9824
rect 8648 9764 8652 9820
rect 8652 9764 8708 9820
rect 8708 9764 8712 9820
rect 8648 9760 8712 9764
rect 8728 9820 8792 9824
rect 8728 9764 8732 9820
rect 8732 9764 8788 9820
rect 8788 9764 8792 9820
rect 8728 9760 8792 9764
rect 8808 9820 8872 9824
rect 8808 9764 8812 9820
rect 8812 9764 8868 9820
rect 8868 9764 8872 9820
rect 8808 9760 8872 9764
rect 60 9692 124 9756
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 7568 9276 7632 9280
rect 7568 9220 7572 9276
rect 7572 9220 7628 9276
rect 7628 9220 7632 9276
rect 7568 9216 7632 9220
rect 7648 9276 7712 9280
rect 7648 9220 7652 9276
rect 7652 9220 7708 9276
rect 7708 9220 7712 9276
rect 7648 9216 7712 9220
rect 7728 9276 7792 9280
rect 7728 9220 7732 9276
rect 7732 9220 7788 9276
rect 7788 9220 7792 9276
rect 7728 9216 7792 9220
rect 7808 9276 7872 9280
rect 7808 9220 7812 9276
rect 7812 9220 7868 9276
rect 7868 9220 7872 9276
rect 7808 9216 7872 9220
rect 8340 9012 8404 9076
rect 3568 8732 3632 8736
rect 3568 8676 3572 8732
rect 3572 8676 3628 8732
rect 3628 8676 3632 8732
rect 3568 8672 3632 8676
rect 3648 8732 3712 8736
rect 3648 8676 3652 8732
rect 3652 8676 3708 8732
rect 3708 8676 3712 8732
rect 3648 8672 3712 8676
rect 3728 8732 3792 8736
rect 3728 8676 3732 8732
rect 3732 8676 3788 8732
rect 3788 8676 3792 8732
rect 3728 8672 3792 8676
rect 3808 8732 3872 8736
rect 3808 8676 3812 8732
rect 3812 8676 3868 8732
rect 3868 8676 3872 8732
rect 3808 8672 3872 8676
rect 8568 8732 8632 8736
rect 8568 8676 8572 8732
rect 8572 8676 8628 8732
rect 8628 8676 8632 8732
rect 8568 8672 8632 8676
rect 8648 8732 8712 8736
rect 8648 8676 8652 8732
rect 8652 8676 8708 8732
rect 8708 8676 8712 8732
rect 8648 8672 8712 8676
rect 8728 8732 8792 8736
rect 8728 8676 8732 8732
rect 8732 8676 8788 8732
rect 8788 8676 8792 8732
rect 8728 8672 8792 8676
rect 8808 8732 8872 8736
rect 8808 8676 8812 8732
rect 8812 8676 8868 8732
rect 8868 8676 8872 8732
rect 8808 8672 8872 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 7568 8188 7632 8192
rect 7568 8132 7572 8188
rect 7572 8132 7628 8188
rect 7628 8132 7632 8188
rect 7568 8128 7632 8132
rect 7648 8188 7712 8192
rect 7648 8132 7652 8188
rect 7652 8132 7708 8188
rect 7708 8132 7712 8188
rect 7648 8128 7712 8132
rect 7728 8188 7792 8192
rect 7728 8132 7732 8188
rect 7732 8132 7788 8188
rect 7788 8132 7792 8188
rect 7728 8128 7792 8132
rect 7808 8188 7872 8192
rect 7808 8132 7812 8188
rect 7812 8132 7868 8188
rect 7868 8132 7872 8188
rect 7808 8128 7872 8132
rect 4108 8060 4172 8124
rect 3568 7644 3632 7648
rect 3568 7588 3572 7644
rect 3572 7588 3628 7644
rect 3628 7588 3632 7644
rect 3568 7584 3632 7588
rect 3648 7644 3712 7648
rect 3648 7588 3652 7644
rect 3652 7588 3708 7644
rect 3708 7588 3712 7644
rect 3648 7584 3712 7588
rect 3728 7644 3792 7648
rect 3728 7588 3732 7644
rect 3732 7588 3788 7644
rect 3788 7588 3792 7644
rect 3728 7584 3792 7588
rect 3808 7644 3872 7648
rect 3808 7588 3812 7644
rect 3812 7588 3868 7644
rect 3868 7588 3872 7644
rect 3808 7584 3872 7588
rect 8568 7644 8632 7648
rect 8568 7588 8572 7644
rect 8572 7588 8628 7644
rect 8628 7588 8632 7644
rect 8568 7584 8632 7588
rect 8648 7644 8712 7648
rect 8648 7588 8652 7644
rect 8652 7588 8708 7644
rect 8708 7588 8712 7644
rect 8648 7584 8712 7588
rect 8728 7644 8792 7648
rect 8728 7588 8732 7644
rect 8732 7588 8788 7644
rect 8788 7588 8792 7644
rect 8728 7584 8792 7588
rect 8808 7644 8872 7648
rect 8808 7588 8812 7644
rect 8812 7588 8868 7644
rect 8868 7588 8872 7644
rect 8808 7584 8872 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 7568 7100 7632 7104
rect 7568 7044 7572 7100
rect 7572 7044 7628 7100
rect 7628 7044 7632 7100
rect 7568 7040 7632 7044
rect 7648 7100 7712 7104
rect 7648 7044 7652 7100
rect 7652 7044 7708 7100
rect 7708 7044 7712 7100
rect 7648 7040 7712 7044
rect 7728 7100 7792 7104
rect 7728 7044 7732 7100
rect 7732 7044 7788 7100
rect 7788 7044 7792 7100
rect 7728 7040 7792 7044
rect 7808 7100 7872 7104
rect 7808 7044 7812 7100
rect 7812 7044 7868 7100
rect 7868 7044 7872 7100
rect 7808 7040 7872 7044
rect 3568 6556 3632 6560
rect 3568 6500 3572 6556
rect 3572 6500 3628 6556
rect 3628 6500 3632 6556
rect 3568 6496 3632 6500
rect 3648 6556 3712 6560
rect 3648 6500 3652 6556
rect 3652 6500 3708 6556
rect 3708 6500 3712 6556
rect 3648 6496 3712 6500
rect 3728 6556 3792 6560
rect 3728 6500 3732 6556
rect 3732 6500 3788 6556
rect 3788 6500 3792 6556
rect 3728 6496 3792 6500
rect 3808 6556 3872 6560
rect 3808 6500 3812 6556
rect 3812 6500 3868 6556
rect 3868 6500 3872 6556
rect 3808 6496 3872 6500
rect 8568 6556 8632 6560
rect 8568 6500 8572 6556
rect 8572 6500 8628 6556
rect 8628 6500 8632 6556
rect 8568 6496 8632 6500
rect 8648 6556 8712 6560
rect 8648 6500 8652 6556
rect 8652 6500 8708 6556
rect 8708 6500 8712 6556
rect 8648 6496 8712 6500
rect 8728 6556 8792 6560
rect 8728 6500 8732 6556
rect 8732 6500 8788 6556
rect 8788 6500 8792 6556
rect 8728 6496 8792 6500
rect 8808 6556 8872 6560
rect 8808 6500 8812 6556
rect 8812 6500 8868 6556
rect 8868 6500 8872 6556
rect 8808 6496 8872 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 7568 6012 7632 6016
rect 7568 5956 7572 6012
rect 7572 5956 7628 6012
rect 7628 5956 7632 6012
rect 7568 5952 7632 5956
rect 7648 6012 7712 6016
rect 7648 5956 7652 6012
rect 7652 5956 7708 6012
rect 7708 5956 7712 6012
rect 7648 5952 7712 5956
rect 7728 6012 7792 6016
rect 7728 5956 7732 6012
rect 7732 5956 7788 6012
rect 7788 5956 7792 6012
rect 7728 5952 7792 5956
rect 7808 6012 7872 6016
rect 7808 5956 7812 6012
rect 7812 5956 7868 6012
rect 7868 5956 7872 6012
rect 7808 5952 7872 5956
rect 3568 5468 3632 5472
rect 3568 5412 3572 5468
rect 3572 5412 3628 5468
rect 3628 5412 3632 5468
rect 3568 5408 3632 5412
rect 3648 5468 3712 5472
rect 3648 5412 3652 5468
rect 3652 5412 3708 5468
rect 3708 5412 3712 5468
rect 3648 5408 3712 5412
rect 3728 5468 3792 5472
rect 3728 5412 3732 5468
rect 3732 5412 3788 5468
rect 3788 5412 3792 5468
rect 3728 5408 3792 5412
rect 3808 5468 3872 5472
rect 3808 5412 3812 5468
rect 3812 5412 3868 5468
rect 3868 5412 3872 5468
rect 3808 5408 3872 5412
rect 8568 5468 8632 5472
rect 8568 5412 8572 5468
rect 8572 5412 8628 5468
rect 8628 5412 8632 5468
rect 8568 5408 8632 5412
rect 8648 5468 8712 5472
rect 8648 5412 8652 5468
rect 8652 5412 8708 5468
rect 8708 5412 8712 5468
rect 8648 5408 8712 5412
rect 8728 5468 8792 5472
rect 8728 5412 8732 5468
rect 8732 5412 8788 5468
rect 8788 5412 8792 5468
rect 8728 5408 8792 5412
rect 8808 5468 8872 5472
rect 8808 5412 8812 5468
rect 8812 5412 8868 5468
rect 8868 5412 8872 5468
rect 8808 5408 8872 5412
rect 7568 4924 7632 4928
rect 7568 4868 7572 4924
rect 7572 4868 7628 4924
rect 7628 4868 7632 4924
rect 7568 4864 7632 4868
rect 7648 4924 7712 4928
rect 7648 4868 7652 4924
rect 7652 4868 7708 4924
rect 7708 4868 7712 4924
rect 7648 4864 7712 4868
rect 7728 4924 7792 4928
rect 7728 4868 7732 4924
rect 7732 4868 7788 4924
rect 7788 4868 7792 4924
rect 7728 4864 7792 4868
rect 7808 4924 7872 4928
rect 7808 4868 7812 4924
rect 7812 4868 7868 4924
rect 7868 4868 7872 4924
rect 7808 4864 7872 4868
rect 1348 4660 1412 4724
rect 3568 4380 3632 4384
rect 3568 4324 3572 4380
rect 3572 4324 3628 4380
rect 3628 4324 3632 4380
rect 3568 4320 3632 4324
rect 3648 4380 3712 4384
rect 3648 4324 3652 4380
rect 3652 4324 3708 4380
rect 3708 4324 3712 4380
rect 3648 4320 3712 4324
rect 3728 4380 3792 4384
rect 3728 4324 3732 4380
rect 3732 4324 3788 4380
rect 3788 4324 3792 4380
rect 3728 4320 3792 4324
rect 3808 4380 3872 4384
rect 3808 4324 3812 4380
rect 3812 4324 3868 4380
rect 3868 4324 3872 4380
rect 3808 4320 3872 4324
rect 8568 4380 8632 4384
rect 8568 4324 8572 4380
rect 8572 4324 8628 4380
rect 8628 4324 8632 4380
rect 8568 4320 8632 4324
rect 8648 4380 8712 4384
rect 8648 4324 8652 4380
rect 8652 4324 8708 4380
rect 8708 4324 8712 4380
rect 8648 4320 8712 4324
rect 8728 4380 8792 4384
rect 8728 4324 8732 4380
rect 8732 4324 8788 4380
rect 8788 4324 8792 4380
rect 8728 4320 8792 4324
rect 8808 4380 8872 4384
rect 8808 4324 8812 4380
rect 8812 4324 8868 4380
rect 8868 4324 8872 4380
rect 8808 4320 8872 4324
rect 7568 3836 7632 3840
rect 7568 3780 7572 3836
rect 7572 3780 7628 3836
rect 7628 3780 7632 3836
rect 7568 3776 7632 3780
rect 7648 3836 7712 3840
rect 7648 3780 7652 3836
rect 7652 3780 7708 3836
rect 7708 3780 7712 3836
rect 7648 3776 7712 3780
rect 7728 3836 7792 3840
rect 7728 3780 7732 3836
rect 7732 3780 7788 3836
rect 7788 3780 7792 3836
rect 7728 3776 7792 3780
rect 7808 3836 7872 3840
rect 7808 3780 7812 3836
rect 7812 3780 7868 3836
rect 7868 3780 7872 3836
rect 7808 3776 7872 3780
rect 3568 3292 3632 3296
rect 3568 3236 3572 3292
rect 3572 3236 3628 3292
rect 3628 3236 3632 3292
rect 3568 3232 3632 3236
rect 3648 3292 3712 3296
rect 3648 3236 3652 3292
rect 3652 3236 3708 3292
rect 3708 3236 3712 3292
rect 3648 3232 3712 3236
rect 3728 3292 3792 3296
rect 3728 3236 3732 3292
rect 3732 3236 3788 3292
rect 3788 3236 3792 3292
rect 3728 3232 3792 3236
rect 3808 3292 3872 3296
rect 3808 3236 3812 3292
rect 3812 3236 3868 3292
rect 3868 3236 3872 3292
rect 3808 3232 3872 3236
rect 8568 3292 8632 3296
rect 8568 3236 8572 3292
rect 8572 3236 8628 3292
rect 8628 3236 8632 3292
rect 8568 3232 8632 3236
rect 8648 3292 8712 3296
rect 8648 3236 8652 3292
rect 8652 3236 8708 3292
rect 8708 3236 8712 3292
rect 8648 3232 8712 3236
rect 8728 3292 8792 3296
rect 8728 3236 8732 3292
rect 8732 3236 8788 3292
rect 8788 3236 8792 3292
rect 8728 3232 8792 3236
rect 8808 3292 8872 3296
rect 8808 3236 8812 3292
rect 8812 3236 8868 3292
rect 8868 3236 8872 3292
rect 8808 3232 8872 3236
rect 4108 2680 4172 2684
rect 4108 2624 4122 2680
rect 4122 2624 4172 2680
rect 4108 2620 4172 2624
rect 7568 2748 7632 2752
rect 7568 2692 7572 2748
rect 7572 2692 7628 2748
rect 7628 2692 7632 2748
rect 7568 2688 7632 2692
rect 7648 2748 7712 2752
rect 7648 2692 7652 2748
rect 7652 2692 7708 2748
rect 7708 2692 7712 2748
rect 7648 2688 7712 2692
rect 7728 2748 7792 2752
rect 7728 2692 7732 2748
rect 7732 2692 7788 2748
rect 7788 2692 7792 2748
rect 7728 2688 7792 2692
rect 7808 2748 7872 2752
rect 7808 2692 7812 2748
rect 7812 2692 7868 2748
rect 7868 2692 7872 2748
rect 7808 2688 7872 2692
rect 8340 2484 8404 2548
rect 3568 2204 3632 2208
rect 3568 2148 3572 2204
rect 3572 2148 3628 2204
rect 3628 2148 3632 2204
rect 3568 2144 3632 2148
rect 3648 2204 3712 2208
rect 3648 2148 3652 2204
rect 3652 2148 3708 2204
rect 3708 2148 3712 2204
rect 3648 2144 3712 2148
rect 3728 2204 3792 2208
rect 3728 2148 3732 2204
rect 3732 2148 3788 2204
rect 3788 2148 3792 2204
rect 3728 2144 3792 2148
rect 3808 2204 3872 2208
rect 3808 2148 3812 2204
rect 3812 2148 3868 2204
rect 3868 2148 3872 2204
rect 3808 2144 3872 2148
rect 8568 2204 8632 2208
rect 8568 2148 8572 2204
rect 8572 2148 8628 2204
rect 8628 2148 8632 2204
rect 8568 2144 8632 2148
rect 8648 2204 8712 2208
rect 8648 2148 8652 2204
rect 8652 2148 8708 2204
rect 8708 2148 8712 2204
rect 8648 2144 8712 2148
rect 8728 2204 8792 2208
rect 8728 2148 8732 2204
rect 8732 2148 8788 2204
rect 8788 2148 8792 2204
rect 8728 2144 8792 2148
rect 8808 2204 8872 2208
rect 8808 2148 8812 2204
rect 8812 2148 8868 2204
rect 8868 2148 8872 2204
rect 8808 2144 8872 2148
rect 7568 1660 7632 1664
rect 7568 1604 7572 1660
rect 7572 1604 7628 1660
rect 7628 1604 7632 1660
rect 7568 1600 7632 1604
rect 7648 1660 7712 1664
rect 7648 1604 7652 1660
rect 7652 1604 7708 1660
rect 7708 1604 7712 1660
rect 7648 1600 7712 1604
rect 7728 1660 7792 1664
rect 7728 1604 7732 1660
rect 7732 1604 7788 1660
rect 7788 1604 7792 1660
rect 7728 1600 7792 1604
rect 7808 1660 7872 1664
rect 7808 1604 7812 1660
rect 7812 1604 7868 1660
rect 7868 1604 7872 1660
rect 7808 1600 7872 1604
rect 60 1592 124 1596
rect 60 1536 110 1592
rect 110 1536 124 1592
rect 60 1532 124 1536
rect 3568 1116 3632 1120
rect 3568 1060 3572 1116
rect 3572 1060 3628 1116
rect 3628 1060 3632 1116
rect 3568 1056 3632 1060
rect 3648 1116 3712 1120
rect 3648 1060 3652 1116
rect 3652 1060 3708 1116
rect 3708 1060 3712 1116
rect 3648 1056 3712 1060
rect 3728 1116 3792 1120
rect 3728 1060 3732 1116
rect 3732 1060 3788 1116
rect 3788 1060 3792 1116
rect 3728 1056 3792 1060
rect 3808 1116 3872 1120
rect 3808 1060 3812 1116
rect 3812 1060 3868 1116
rect 3868 1060 3872 1116
rect 3808 1056 3872 1060
rect 8568 1116 8632 1120
rect 8568 1060 8572 1116
rect 8572 1060 8628 1116
rect 8628 1060 8632 1116
rect 8568 1056 8632 1060
rect 8648 1116 8712 1120
rect 8648 1060 8652 1116
rect 8652 1060 8708 1116
rect 8708 1060 8712 1116
rect 8648 1056 8712 1060
rect 8728 1116 8792 1120
rect 8728 1060 8732 1116
rect 8732 1060 8788 1116
rect 8788 1060 8792 1116
rect 8728 1056 8792 1060
rect 8808 1116 8872 1120
rect 8808 1060 8812 1116
rect 8812 1060 8868 1116
rect 8868 1060 8872 1116
rect 8808 1056 8872 1060
<< metal4 >>
rect 2560 15808 2880 15824
rect 2560 15744 2568 15808
rect 2632 15744 2648 15808
rect 2712 15744 2728 15808
rect 2792 15744 2808 15808
rect 2872 15744 2880 15808
rect 979 15332 1045 15333
rect 979 15268 980 15332
rect 1044 15268 1045 15332
rect 979 15267 1045 15268
rect 982 12477 1042 15267
rect 2560 14720 2880 15744
rect 2560 14656 2568 14720
rect 2632 14656 2648 14720
rect 2712 14656 2728 14720
rect 2792 14656 2808 14720
rect 2872 14656 2880 14720
rect 2560 13632 2880 14656
rect 2560 13568 2568 13632
rect 2632 13568 2648 13632
rect 2712 13568 2728 13632
rect 2792 13568 2808 13632
rect 2872 13568 2880 13632
rect 2560 13206 2880 13568
rect 2560 12970 2602 13206
rect 2838 12970 2880 13206
rect 2560 12544 2880 12970
rect 2560 12480 2568 12544
rect 2632 12480 2648 12544
rect 2712 12480 2728 12544
rect 2792 12480 2808 12544
rect 2872 12480 2880 12544
rect 979 12476 1045 12477
rect 979 12412 980 12476
rect 1044 12412 1045 12476
rect 979 12411 1045 12412
rect 1347 12476 1413 12477
rect 1347 12412 1348 12476
rect 1412 12412 1413 12476
rect 1347 12411 1413 12412
rect 59 9756 125 9757
rect 59 9692 60 9756
rect 124 9692 125 9756
rect 59 9691 125 9692
rect 62 1597 122 9691
rect 1350 4725 1410 12411
rect 2560 11456 2880 12480
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9206 2880 9216
rect 2560 8970 2602 9206
rect 2838 8970 2880 9206
rect 2560 8192 2880 8970
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 7104 2880 8128
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5206 2880 5952
rect 2560 4970 2602 5206
rect 2838 4970 2880 5206
rect 2560 4893 2880 4970
rect 3560 15264 3880 15824
rect 3560 15200 3568 15264
rect 3632 15200 3648 15264
rect 3712 15200 3728 15264
rect 3792 15200 3808 15264
rect 3872 15200 3880 15264
rect 3560 14206 3880 15200
rect 3560 14176 3602 14206
rect 3838 14176 3880 14206
rect 3560 14112 3568 14176
rect 3872 14112 3880 14176
rect 3560 13970 3602 14112
rect 3838 13970 3880 14112
rect 3560 13088 3880 13970
rect 3560 13024 3568 13088
rect 3632 13024 3648 13088
rect 3712 13024 3728 13088
rect 3792 13024 3808 13088
rect 3872 13024 3880 13088
rect 3560 12000 3880 13024
rect 3560 11936 3568 12000
rect 3632 11936 3648 12000
rect 3712 11936 3728 12000
rect 3792 11936 3808 12000
rect 3872 11936 3880 12000
rect 3560 10912 3880 11936
rect 3560 10848 3568 10912
rect 3632 10848 3648 10912
rect 3712 10848 3728 10912
rect 3792 10848 3808 10912
rect 3872 10848 3880 10912
rect 3560 10206 3880 10848
rect 3560 9970 3602 10206
rect 3838 9970 3880 10206
rect 3560 9824 3880 9970
rect 3560 9760 3568 9824
rect 3632 9760 3648 9824
rect 3712 9760 3728 9824
rect 3792 9760 3808 9824
rect 3872 9760 3880 9824
rect 3560 8736 3880 9760
rect 3560 8672 3568 8736
rect 3632 8672 3648 8736
rect 3712 8672 3728 8736
rect 3792 8672 3808 8736
rect 3872 8672 3880 8736
rect 3560 7648 3880 8672
rect 4560 15206 4880 15824
rect 4560 14970 4602 15206
rect 4838 14970 4880 15206
rect 4560 11206 4880 14970
rect 4560 10970 4602 11206
rect 4838 10970 4880 11206
rect 4107 8124 4173 8125
rect 4107 8060 4108 8124
rect 4172 8060 4173 8124
rect 4107 8059 4173 8060
rect 3560 7584 3568 7648
rect 3632 7584 3648 7648
rect 3712 7584 3728 7648
rect 3792 7584 3808 7648
rect 3872 7584 3880 7648
rect 3560 6560 3880 7584
rect 3560 6496 3568 6560
rect 3632 6496 3648 6560
rect 3712 6496 3728 6560
rect 3792 6496 3808 6560
rect 3872 6496 3880 6560
rect 3560 6206 3880 6496
rect 3560 5970 3602 6206
rect 3838 5970 3880 6206
rect 3560 5472 3880 5970
rect 3560 5408 3568 5472
rect 3632 5408 3648 5472
rect 3712 5408 3728 5472
rect 3792 5408 3808 5472
rect 3872 5408 3880 5472
rect 1347 4724 1413 4725
rect 1347 4660 1348 4724
rect 1412 4660 1413 4724
rect 1347 4659 1413 4660
rect 3560 4384 3880 5408
rect 3560 4320 3568 4384
rect 3632 4320 3648 4384
rect 3712 4320 3728 4384
rect 3792 4320 3808 4384
rect 3872 4320 3880 4384
rect 1996 4206 2276 4248
rect 1996 3970 2018 4206
rect 2254 3970 2276 4206
rect 1996 3928 2276 3970
rect 3560 3296 3880 4320
rect 1256 3206 1536 3248
rect 1256 2970 1278 3206
rect 1514 2970 1536 3206
rect 1256 2928 1536 2970
rect 3560 3232 3568 3296
rect 3632 3232 3648 3296
rect 3712 3232 3728 3296
rect 3792 3232 3808 3296
rect 3872 3232 3880 3296
rect 3560 2208 3880 3232
rect 4110 2685 4170 8059
rect 4560 7206 4880 10970
rect 4560 6970 4602 7206
rect 4838 6970 4880 7206
rect 4560 3206 4880 6970
rect 4560 2970 4602 3206
rect 4838 2970 4880 3206
rect 4107 2684 4173 2685
rect 4107 2620 4108 2684
rect 4172 2620 4173 2684
rect 4107 2619 4173 2620
rect 3560 2144 3568 2208
rect 3632 2206 3648 2208
rect 3712 2206 3728 2208
rect 3792 2206 3808 2208
rect 3872 2144 3880 2208
rect 3560 1970 3602 2144
rect 3838 1970 3880 2144
rect 59 1596 125 1597
rect 59 1532 60 1596
rect 124 1532 125 1596
rect 59 1531 125 1532
rect 3560 1120 3880 1970
rect 3560 1056 3568 1120
rect 3632 1056 3648 1120
rect 3712 1056 3728 1120
rect 3792 1056 3808 1120
rect 3872 1056 3880 1120
rect 3560 1040 3880 1056
rect 4560 1040 4880 2970
rect 5560 4206 5880 15824
rect 5560 3970 5602 4206
rect 5838 3970 5880 4206
rect 5560 1040 5880 3970
rect 7560 15808 7880 15824
rect 7560 15744 7568 15808
rect 7632 15744 7648 15808
rect 7712 15744 7728 15808
rect 7792 15744 7808 15808
rect 7872 15744 7880 15808
rect 7560 14720 7880 15744
rect 7560 14656 7568 14720
rect 7632 14656 7648 14720
rect 7712 14656 7728 14720
rect 7792 14656 7808 14720
rect 7872 14656 7880 14720
rect 7560 13632 7880 14656
rect 7560 13568 7568 13632
rect 7632 13568 7648 13632
rect 7712 13568 7728 13632
rect 7792 13568 7808 13632
rect 7872 13568 7880 13632
rect 7560 13206 7880 13568
rect 7560 12970 7602 13206
rect 7838 12970 7880 13206
rect 7560 12544 7880 12970
rect 8560 15264 8880 15824
rect 8560 15200 8568 15264
rect 8632 15200 8648 15264
rect 8712 15200 8728 15264
rect 8792 15200 8808 15264
rect 8872 15200 8880 15264
rect 8560 14206 8880 15200
rect 8560 14176 8602 14206
rect 8838 14176 8880 14206
rect 8560 14112 8568 14176
rect 8872 14112 8880 14176
rect 8560 13970 8602 14112
rect 8838 13970 8880 14112
rect 8560 13088 8880 13970
rect 8560 13024 8568 13088
rect 8632 13024 8648 13088
rect 8712 13024 8728 13088
rect 8792 13024 8808 13088
rect 8872 13024 8880 13088
rect 7971 12884 8037 12885
rect 7971 12820 7972 12884
rect 8036 12820 8037 12884
rect 7971 12819 8037 12820
rect 7974 12613 8034 12819
rect 7971 12612 8037 12613
rect 7971 12548 7972 12612
rect 8036 12548 8037 12612
rect 7971 12547 8037 12548
rect 7560 12480 7568 12544
rect 7632 12480 7648 12544
rect 7712 12480 7728 12544
rect 7792 12480 7808 12544
rect 7872 12480 7880 12544
rect 7560 11456 7880 12480
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 7560 10368 7880 11392
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 9280 7880 10304
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 9206 7880 9216
rect 7560 8970 7602 9206
rect 7838 8970 7880 9206
rect 8560 12000 8880 13024
rect 8560 11936 8568 12000
rect 8632 11936 8648 12000
rect 8712 11936 8728 12000
rect 8792 11936 8808 12000
rect 8872 11936 8880 12000
rect 8560 10912 8880 11936
rect 8560 10848 8568 10912
rect 8632 10848 8648 10912
rect 8712 10848 8728 10912
rect 8792 10848 8808 10912
rect 8872 10848 8880 10912
rect 8560 10206 8880 10848
rect 8560 9970 8602 10206
rect 8838 9970 8880 10206
rect 8560 9824 8880 9970
rect 8560 9760 8568 9824
rect 8632 9760 8648 9824
rect 8712 9760 8728 9824
rect 8792 9760 8808 9824
rect 8872 9760 8880 9824
rect 8339 9076 8405 9077
rect 8339 9012 8340 9076
rect 8404 9012 8405 9076
rect 8339 9011 8405 9012
rect 7560 8192 7880 8970
rect 7560 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7880 8192
rect 7560 7104 7880 8128
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 6016 7880 7040
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 5206 7880 5952
rect 7560 4970 7602 5206
rect 7838 4970 7880 5206
rect 7560 4928 7880 4970
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 7560 3840 7880 4864
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 2752 7880 3776
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 1664 7880 2688
rect 8342 2549 8402 9011
rect 8560 8736 8880 9760
rect 8560 8672 8568 8736
rect 8632 8672 8648 8736
rect 8712 8672 8728 8736
rect 8792 8672 8808 8736
rect 8872 8672 8880 8736
rect 8560 7648 8880 8672
rect 8560 7584 8568 7648
rect 8632 7584 8648 7648
rect 8712 7584 8728 7648
rect 8792 7584 8808 7648
rect 8872 7584 8880 7648
rect 8560 6560 8880 7584
rect 8560 6496 8568 6560
rect 8632 6496 8648 6560
rect 8712 6496 8728 6560
rect 8792 6496 8808 6560
rect 8872 6496 8880 6560
rect 8560 6206 8880 6496
rect 8560 5970 8602 6206
rect 8838 5970 8880 6206
rect 8560 5472 8880 5970
rect 8560 5408 8568 5472
rect 8632 5408 8648 5472
rect 8712 5408 8728 5472
rect 8792 5408 8808 5472
rect 8872 5408 8880 5472
rect 8560 4384 8880 5408
rect 8560 4320 8568 4384
rect 8632 4320 8648 4384
rect 8712 4320 8728 4384
rect 8792 4320 8808 4384
rect 8872 4320 8880 4384
rect 8560 3296 8880 4320
rect 8560 3232 8568 3296
rect 8632 3232 8648 3296
rect 8712 3232 8728 3296
rect 8792 3232 8808 3296
rect 8872 3232 8880 3296
rect 8339 2548 8405 2549
rect 8339 2484 8340 2548
rect 8404 2484 8405 2548
rect 8339 2483 8405 2484
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 7560 1206 7880 1600
rect 7560 970 7602 1206
rect 7838 970 7880 1206
rect 8560 2208 8880 3232
rect 8560 2144 8568 2208
rect 8632 2206 8648 2208
rect 8712 2206 8728 2208
rect 8792 2206 8808 2208
rect 8872 2144 8880 2208
rect 8560 1970 8602 2144
rect 8838 1970 8880 2144
rect 8560 1120 8880 1970
rect 8560 1056 8568 1120
rect 8632 1056 8648 1120
rect 8712 1056 8728 1120
rect 8792 1056 8808 1120
rect 8872 1056 8880 1120
rect 8560 1040 8880 1056
rect 9560 15206 9880 15824
rect 9560 14970 9602 15206
rect 9838 14970 9880 15206
rect 9560 11206 9880 14970
rect 9560 10970 9602 11206
rect 9838 10970 9880 11206
rect 9560 7206 9880 10970
rect 9560 6970 9602 7206
rect 9838 6970 9880 7206
rect 9560 3206 9880 6970
rect 9560 2970 9602 3206
rect 9838 2970 9880 3206
rect 9560 1040 9880 2970
rect 7560 928 7880 970
<< via4 >>
rect 2602 12970 2838 13206
rect 2602 8970 2838 9206
rect 2602 4970 2838 5206
rect 3602 14176 3838 14206
rect 3602 14112 3632 14176
rect 3632 14112 3648 14176
rect 3648 14112 3712 14176
rect 3712 14112 3728 14176
rect 3728 14112 3792 14176
rect 3792 14112 3808 14176
rect 3808 14112 3838 14176
rect 3602 13970 3838 14112
rect 3602 9970 3838 10206
rect 4602 14970 4838 15206
rect 4602 10970 4838 11206
rect 3602 5970 3838 6206
rect 2018 3970 2254 4206
rect 1278 2970 1514 3206
rect 4602 6970 4838 7206
rect 4602 2970 4838 3206
rect 3602 2144 3632 2206
rect 3632 2144 3648 2206
rect 3648 2144 3712 2206
rect 3712 2144 3728 2206
rect 3728 2144 3792 2206
rect 3792 2144 3808 2206
rect 3808 2144 3838 2206
rect 3602 1970 3838 2144
rect 5602 3970 5838 4206
rect 7602 12970 7838 13206
rect 8602 14176 8838 14206
rect 8602 14112 8632 14176
rect 8632 14112 8648 14176
rect 8648 14112 8712 14176
rect 8712 14112 8728 14176
rect 8728 14112 8792 14176
rect 8792 14112 8808 14176
rect 8808 14112 8838 14176
rect 8602 13970 8838 14112
rect 7602 8970 7838 9206
rect 8602 9970 8838 10206
rect 7602 4970 7838 5206
rect 8602 5970 8838 6206
rect 7602 970 7838 1206
rect 8602 2144 8632 2206
rect 8632 2144 8648 2206
rect 8648 2144 8712 2206
rect 8712 2144 8728 2206
rect 8728 2144 8792 2206
rect 8792 2144 8808 2206
rect 8808 2144 8838 2206
rect 8602 1970 8838 2144
rect 9602 14970 9838 15206
rect 9602 10970 9838 11206
rect 9602 6970 9838 7206
rect 9602 2970 9838 3206
<< metal5 >>
rect 872 15206 9892 15248
rect 872 14970 4602 15206
rect 4838 14970 9602 15206
rect 9838 14970 9892 15206
rect 872 14928 9892 14970
rect 872 14206 9892 14248
rect 872 13970 3602 14206
rect 3838 13970 8602 14206
rect 8838 13970 9892 14206
rect 872 13928 9892 13970
rect 872 13206 9892 13248
rect 872 12970 2602 13206
rect 2838 12970 7602 13206
rect 7838 12970 9892 13206
rect 872 12928 9892 12970
rect 872 11206 9892 11248
rect 872 10970 4602 11206
rect 4838 10970 9602 11206
rect 9838 10970 9892 11206
rect 872 10928 9892 10970
rect 872 10206 9892 10248
rect 872 9970 3602 10206
rect 3838 9970 8602 10206
rect 8838 9970 9892 10206
rect 872 9928 9892 9970
rect 872 9206 9892 9248
rect 872 8970 2602 9206
rect 2838 8970 7602 9206
rect 7838 8970 9892 9206
rect 872 8928 9892 8970
rect 872 7206 9892 7248
rect 872 6970 4602 7206
rect 4838 6970 9602 7206
rect 9838 6970 9892 7206
rect 872 6928 9892 6970
rect 872 6206 9892 6248
rect 872 5970 3602 6206
rect 3838 5970 8602 6206
rect 8838 5970 9892 6206
rect 872 5928 9892 5970
rect 872 5206 9892 5248
rect 872 4970 2602 5206
rect 2838 4970 7602 5206
rect 7838 4970 9892 5206
rect 872 4928 9892 4970
rect 872 4206 9892 4248
rect 872 3970 2018 4206
rect 2254 3970 5602 4206
rect 5838 3970 9892 4206
rect 872 3928 9892 3970
rect 872 3206 9892 3248
rect 872 2970 1278 3206
rect 1514 2970 4602 3206
rect 4838 2970 9602 3206
rect 9838 2970 9892 3206
rect 872 2928 9892 2970
rect 872 2206 9892 2248
rect 872 1970 3602 2206
rect 3838 1970 8602 2206
rect 8838 1970 9892 2206
rect 872 1928 9892 1970
rect 872 1206 9892 1248
rect 872 970 7602 1206
rect 7838 970 9892 1206
rect 872 928 9892 970
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 0
transform 1 0 3312 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31
timestamp 0
transform 1 0 3772 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 0
transform 1 0 4416 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45
timestamp 0
transform 1 0 5060 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52
timestamp 0
transform 1 0 5704 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 0
transform 1 0 6164 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64
timestamp 0
transform 1 0 6808 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71
timestamp 0
transform 1 0 7452 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80
timestamp 0
transform 1 0 8280 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92
timestamp 0
transform 1 0 9384 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 0
transform 1 0 3312 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_31
timestamp 0
transform 1 0 3772 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 0
transform 1 0 4416 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 0
transform 1 0 5060 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 0
transform 1 0 5704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_59
timestamp 0
transform 1 0 6348 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_66
timestamp 0
transform 1 0 6992 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_73
timestamp 0
transform 1 0 7636 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_80
timestamp 0
transform 1 0 8280 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 0
transform 1 0 8740 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 0
transform 1 0 9384 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_31
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 0
transform 1 0 4508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_44
timestamp 0
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_50
timestamp 0
transform 1 0 5520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_52
timestamp 0
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 0
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_71
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_79
timestamp 0
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 0
transform 1 0 8740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_92
timestamp 0
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 0
transform 1 0 3312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 0
transform 1 0 4324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_44
timestamp 0
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 0
transform 1 0 5612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_58
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 0
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_76
timestamp 0
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_80
timestamp 0
transform 1 0 8280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 0
transform 1 0 8740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 0
transform 1 0 9384 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 0
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_31
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_38
timestamp 0
transform 1 0 4416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_42
timestamp 0
transform 1 0 4784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_46
timestamp 0
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_50
timestamp 0
transform 1 0 5520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_52
timestamp 0
transform 1 0 5704 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_57
timestamp 0
transform 1 0 6164 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_65
timestamp 0
transform 1 0 6900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_69
timestamp 0
transform 1 0 7268 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 0
transform 1 0 8004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_82
timestamp 0
transform 1 0 8464 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_92
timestamp 0
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_26
timestamp 0
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 0
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 0
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 0
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_59
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp 0
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_67
timestamp 0
transform 1 0 7084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_74
timestamp 0
transform 1 0 7728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_78
timestamp 0
transform 1 0 8096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_80
timestamp 0
transform 1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 0
transform 1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 0
transform 1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_31
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 0
transform 1 0 4784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_49
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_52
timestamp 0
transform 1 0 5704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 0
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_65
timestamp 0
transform 1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_72
timestamp 0
transform 1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp 0
transform 1 0 8280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_84
timestamp 0
transform 1 0 8648 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_92
timestamp 0
transform 1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_26
timestamp 0
transform 1 0 3312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_32
timestamp 0
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_36
timestamp 0
transform 1 0 4232 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_44
timestamp 0
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_54
timestamp 0
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_58
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_64
timestamp 0
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_71
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_80
timestamp 0
transform 1 0 8280 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_86
timestamp 0
transform 1 0 8832 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_91
timestamp 0
transform 1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 0
transform 1 0 1196 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 0
transform 1 0 1564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 0
transform 1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 0
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 0
transform 1 0 5612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_55
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_57
timestamp 0
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_67
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_75
timestamp 0
transform 1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 0
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_91
timestamp 0
transform 1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 0
transform 1 0 1196 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 0
transform 1 0 1564 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_16
timestamp 0
transform 1 0 2392 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_24
timestamp 0
transform 1 0 3128 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 0
transform 1 0 5060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_49
timestamp 0
transform 1 0 5428 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 0
transform 1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_87
timestamp 0
transform 1 0 8924 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_93
timestamp 0
transform 1 0 9476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 0
transform 1 0 1196 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 0
transform 1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_52
timestamp 0
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 0
transform 1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_92
timestamp 0
transform 1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 0
transform 1 0 1196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 0
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 0
transform 1 0 3680 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 0
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 0
transform 1 0 8740 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 0
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 0
transform 1 0 1196 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 0
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_39
timestamp 0
transform 1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_67
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 0
transform 1 0 8556 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_92
timestamp 0
transform 1 0 9384 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 0
transform 1 0 1196 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 0
transform 1 0 1564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_16
timestamp 0
transform 1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_46
timestamp 0
transform 1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 0
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_67
timestamp 0
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp 0
transform 1 0 9384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 0
transform 1 0 1196 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 0
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp 0
transform 1 0 3956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_42
timestamp 0
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 0
transform 1 0 5152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_67
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 0
transform 1 0 8004 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 0
transform 1 0 8556 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_91
timestamp 0
transform 1 0 9292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 0
transform 1 0 1196 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 0
transform 1 0 3128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 0
transform 1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 0
transform 1 0 6992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_90
timestamp 0
transform 1 0 9200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 0
transform 1 0 1196 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_14
timestamp 0
transform 1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 0
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_51
timestamp 0
transform 1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 0
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_92
timestamp 0
transform 1 0 9384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 0
transform 1 0 1196 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_10
timestamp 0
transform 1 0 1840 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_16
timestamp 0
transform 1 0 2392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_43
timestamp 0
transform 1 0 4876 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 0
transform 1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 0
transform 1 0 8740 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_92
timestamp 0
transform 1 0 9384 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 0
transform 1 0 1196 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 0
transform 1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 0
transform 1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_29
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_35
timestamp 0
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_44
timestamp 0
transform 1 0 4968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_48
timestamp 0
transform 1 0 5336 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 0
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 0
transform 1 0 8096 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_91
timestamp 0
transform 1 0 9292 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 0
transform 1 0 1196 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 0
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_30
timestamp 0
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 0
transform 1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_79
timestamp 0
transform 1 0 8188 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_91
timestamp 0
transform 1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 0
transform 1 0 1196 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 0
transform 1 0 3312 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 0
transform 1 0 4048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_64
timestamp 0
transform 1 0 6808 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_70
timestamp 0
transform 1 0 7360 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 0
transform 1 0 8556 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_92
timestamp 0
transform 1 0 9384 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 0
transform 1 0 1196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_14
timestamp 0
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_44
timestamp 0
transform 1 0 4968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 0
transform 1 0 5888 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_81
timestamp 0
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_85
timestamp 0
transform 1 0 8740 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp 0
transform 1 0 9384 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 0
transform 1 0 1196 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 0
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_40
timestamp 0
transform 1 0 4600 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_72
timestamp 0
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_76
timestamp 0
transform 1 0 7912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 0
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_91
timestamp 0
transform 1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 0
transform 1 0 1196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_14
timestamp 0
transform 1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_44
timestamp 0
transform 1 0 4968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_48
timestamp 0
transform 1 0 5336 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 0
transform 1 0 5888 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 0
transform 1 0 6532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_88
timestamp 0
transform 1 0 9016 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 0
transform 1 0 1196 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 0
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_34
timestamp 0
transform 1 0 4048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_43
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_67
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 0
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_92
timestamp 0
transform 1 0 9384 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 0
transform 1 0 1196 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_11
timestamp 0
transform 1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 0
transform 1 0 2300 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 0
transform 1 0 2852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 0
transform 1 0 3680 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_42
timestamp 0
transform 1 0 4784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 0
transform 1 0 5888 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_61
timestamp 0
transform 1 0 6532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_82
timestamp 0
transform 1 0 8464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_86
timestamp 0
transform 1 0 8832 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_91
timestamp 0
transform 1 0 9292 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 0
transform 1 0 1196 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_10
timestamp 0
transform 1 0 1840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_18
timestamp 0
transform 1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 0
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_46
timestamp 0
transform 1 0 5152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_54
timestamp 0
transform 1 0 5888 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_57
timestamp 0
transform 1 0 6164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 0
transform 1 0 6532 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 0
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_91
timestamp 0
transform 1 0 9292 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 920 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 9844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 920 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 9844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 920 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 9844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 920 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 9844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 920 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 920 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 9844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 920 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 9844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 920 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 0
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 0
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 0
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 0
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 0
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 0
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 0
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 0
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 0
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 0
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 0
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 0
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 0
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 0
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 0
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 0
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 0
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 0
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 0
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 0
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 0
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 0
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 0
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 0
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 0
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 0
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 0
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 0
transform 1 0 6072 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 0
transform 1 0 3496 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 0
transform 1 0 8648 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 0
transform 1 0 6072 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 0
transform 1 0 3496 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 0
transform 1 0 8648 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 0
transform 1 0 6072 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 0
transform 1 0 3496 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 0
transform 1 0 8648 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 0
transform 1 0 6072 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 0
transform 1 0 3496 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 0
transform 1 0 6072 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 0
transform 1 0 8648 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _085_
timestamp 0
transform 1 0 6440 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _086_
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _087_
timestamp 0
transform -1 0 6808 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _088_
timestamp 0
transform -1 0 9384 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _089_
timestamp 0
transform -1 0 9292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _090_
timestamp 0
transform 1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _091_
timestamp 0
transform -1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _093_
timestamp 0
transform -1 0 6992 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _094_
timestamp 0
transform 1 0 8924 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _095_
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 0
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _097_
timestamp 0
transform -1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _098_
timestamp 0
transform 1 0 2944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _099_
timestamp 0
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _100_
timestamp 0
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 0
transform -1 0 9384 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _102_
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _103_
timestamp 0
transform 1 0 2392 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 0
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _105_
timestamp 0
transform 1 0 5336 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _106__5
timestamp 0
transform -1 0 6164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp 0
transform -1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _108_
timestamp 0
transform 1 0 7452 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _109_
timestamp 0
transform 1 0 4784 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _110_
timestamp 0
transform 1 0 1472 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 0
transform -1 0 4416 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112__6
timestamp 0
transform -1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _113_
timestamp 0
transform 1 0 6072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _114_
timestamp 0
transform 1 0 4416 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 0
transform -1 0 4784 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116__7
timestamp 0
transform 1 0 3496 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _117_
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _118_
timestamp 0
transform -1 0 5888 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 0
transform -1 0 5704 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120__8
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _121_
timestamp 0
transform 1 0 6072 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 0
transform 1 0 7636 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 0
transform -1 0 3772 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124__9
timestamp 0
transform -1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _125_
timestamp 0
transform 1 0 5888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _126_
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 0
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _128__10
timestamp 0
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _129_
timestamp 0
transform 1 0 3496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _130_
timestamp 0
transform 1 0 3220 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 0
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _132__11
timestamp 0
transform 1 0 7360 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _133_
timestamp 0
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _134_
timestamp 0
transform 1 0 5428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 0
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136__12
timestamp 0
transform -1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _137_
timestamp 0
transform -1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _138_
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 0
transform -1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _140__13
timestamp 0
transform 1 0 9108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _141_
timestamp 0
transform 1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _142_
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 0
transform -1 0 6256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144__14
timestamp 0
transform 1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _145_
timestamp 0
transform 1 0 6992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _146_
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 0
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148__1
timestamp 0
transform -1 0 4232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _149_
timestamp 0
transform 1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _150_
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 0
transform -1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _152__2
timestamp 0
transform -1 0 6900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _153_
timestamp 0
transform 1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _154_
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 0
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156__3
timestamp 0
transform 1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _157_
timestamp 0
transform 1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _158__4
timestamp 0
transform 1 0 4784 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _159_
timestamp 0
transform -1 0 4968 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _160_
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _161_
timestamp 0
transform 1 0 4416 0 1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _162_
timestamp 0
transform 1 0 5152 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _163_
timestamp 0
transform 1 0 2760 0 -1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _164_
timestamp 0
transform 1 0 3496 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _165_
timestamp 0
transform 1 0 2576 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _166_
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _167_
timestamp 0
transform -1 0 8740 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _168_
timestamp 0
transform -1 0 9016 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _169_
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _170_
timestamp 0
transform 1 0 6072 0 1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _171_
timestamp 0
transform 1 0 6532 0 -1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__dfrtp_1  _172_
timestamp 0
transform -1 0 8464 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _173_
timestamp 0
transform -1 0 3312 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _174_
timestamp 0
transform -1 0 3312 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _175_
timestamp 0
transform 1 0 1472 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _176_
timestamp 0
transform 1 0 1472 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _177_
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _178_
timestamp 0
transform -1 0 5704 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _179_
timestamp 0
transform 1 0 4048 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _180_
timestamp 0
transform -1 0 5060 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _181_
timestamp 0
transform -1 0 3680 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _182_
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _183_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _184_
timestamp 0
transform 1 0 6532 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _185_
timestamp 0
transform -1 0 8464 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 0
transform -1 0 4416 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _187_
timestamp 0
transform -1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _188_
timestamp 0
transform -1 0 1840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_8  _189_
timestamp 0
transform -1 0 9384 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__068_
timestamp 0
transform -1 0 5888 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock
timestamp 0
transform -1 0 7268 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 0
transform -1 0 9200 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__068_
timestamp 0
transform 1 0 1472 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_clock
timestamp 0
transform -1 0 3680 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_load
timestamp 0
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__068_
timestamp 0
transform 1 0 1472 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_clock
timestamp 0
transform 1 0 5244 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_load
timestamp 0
transform -1 0 7084 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  const_source
timestamp 0
transform -1 0 8740 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 0
transform -1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 0
transform -1 0 9384 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf
timestamp 0
transform 1 0 1472 0 -1 9792
box -38 -48 1694 592
use gpio_logic_high  gpio_logic_high
timestamp 0
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform 1 0 1472 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform 1 0 1656 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform 1 0 4048 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform 1 0 1656 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform 1 0 7636 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform 1 0 7452 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform 1 0 1472 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform 1 0 4048 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform 1 0 2576 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform 1 0 6348 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform 1 0 5152 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform -1 0 8188 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform -1 0 5888 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 0
transform 1 0 1472 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 0
transform 1 0 1472 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 0
transform -1 0 4968 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 0
transform 1 0 2576 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output1
timestamp 0
transform 1 0 9016 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 0
transform -1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 0
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 0
transform 1 0 9016 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 0
transform -1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 0
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform -1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform 1 0 8924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform -1 0 2760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform 1 0 8004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform 1 0 5520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  output15
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output16
timestamp 0
transform -1 0 5152 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output17
timestamp 0
transform 1 0 3496 0 -1 3264
box -38 -48 866 592
<< labels >>
flabel metal2 s 938 16200 994 17000 0 FreeSans 280 90 0 0 gpio_defaults[0]
port 1 nsew
flabel metal2 s 5538 16200 5594 17000 0 FreeSans 280 90 0 0 gpio_defaults[10]
port 2 nsew
flabel metal2 s 5998 16200 6054 17000 0 FreeSans 280 90 0 0 gpio_defaults[11]
port 3 nsew
flabel metal2 s 6458 16200 6514 17000 0 FreeSans 280 90 0 0 gpio_defaults[12]
port 4 nsew
flabel metal2 s 1398 16200 1454 17000 0 FreeSans 280 90 0 0 gpio_defaults[1]
port 5 nsew
flabel metal2 s 1858 16200 1914 17000 0 FreeSans 280 90 0 0 gpio_defaults[2]
port 6 nsew
flabel metal2 s 2318 16200 2374 17000 0 FreeSans 280 90 0 0 gpio_defaults[3]
port 7 nsew
flabel metal2 s 2778 16200 2834 17000 0 FreeSans 280 90 0 0 gpio_defaults[4]
port 8 nsew
flabel metal2 s 3238 16200 3294 17000 0 FreeSans 280 90 0 0 gpio_defaults[5]
port 9 nsew
flabel metal2 s 3698 16200 3754 17000 0 FreeSans 280 90 0 0 gpio_defaults[6]
port 10 nsew
flabel metal2 s 4158 16200 4214 17000 0 FreeSans 280 90 0 0 gpio_defaults[7]
port 11 nsew
flabel metal2 s 4618 16200 4674 17000 0 FreeSans 280 90 0 0 gpio_defaults[8]
port 12 nsew
flabel metal2 s 5078 16200 5134 17000 0 FreeSans 280 90 0 0 gpio_defaults[9]
port 13 nsew
flabel metal3 s 14000 4904 34000 5024 0 FreeSans 600 0 0 0 mgmt_gpio_in
port 14 nsew
flabel metal3 s 14000 5720 34000 5840 0 FreeSans 600 0 0 0 mgmt_gpio_oeb
port 15 nsew
flabel metal3 s 14000 6128 34000 6248 0 FreeSans 600 0 0 0 mgmt_gpio_out
port 16 nsew
flabel metal3 s 14000 5312 34000 5432 0 FreeSans 600 0 0 0 one
port 17 nsew
flabel metal3 s 14000 6536 34000 6656 0 FreeSans 600 0 0 0 pad_gpio_ana_en
port 18 nsew
flabel metal3 s 14000 6944 34000 7064 0 FreeSans 600 0 0 0 pad_gpio_ana_pol
port 19 nsew
flabel metal3 s 14000 7352 34000 7472 0 FreeSans 600 0 0 0 pad_gpio_ana_sel
port 20 nsew
flabel metal3 s 14000 7760 34000 7880 0 FreeSans 600 0 0 0 pad_gpio_dm[0]
port 21 nsew
flabel metal3 s 14000 8168 34000 8288 0 FreeSans 600 0 0 0 pad_gpio_dm[1]
port 22 nsew
flabel metal3 s 14000 8576 34000 8696 0 FreeSans 600 0 0 0 pad_gpio_dm[2]
port 23 nsew
flabel metal3 s 14000 8984 34000 9104 0 FreeSans 600 0 0 0 pad_gpio_holdover
port 24 nsew
flabel metal3 s 14000 9392 34000 9512 0 FreeSans 600 0 0 0 pad_gpio_ib_mode_sel
port 25 nsew
flabel metal3 s 14000 9800 34000 9920 0 FreeSans 600 0 0 0 pad_gpio_in
port 26 nsew
flabel metal3 s 14000 10208 34000 10328 0 FreeSans 600 0 0 0 pad_gpio_inenb
port 27 nsew
flabel metal3 s 14000 10616 34000 10736 0 FreeSans 600 0 0 0 pad_gpio_out
port 28 nsew
flabel metal3 s 14000 11024 34000 11144 0 FreeSans 600 0 0 0 pad_gpio_outenb
port 29 nsew
flabel metal3 s 14000 11432 34000 11552 0 FreeSans 600 0 0 0 pad_gpio_slow_sel
port 30 nsew
flabel metal3 s 14000 11840 34000 11960 0 FreeSans 600 0 0 0 pad_gpio_vtrip_sel
port 31 nsew
flabel metal3 s 14000 12248 34000 12368 0 FreeSans 600 0 0 0 resetn
port 32 nsew
flabel metal3 s 14000 12656 34000 12776 0 FreeSans 600 0 0 0 resetn_out
port 33 nsew
flabel metal3 s 14000 13064 34000 13184 0 FreeSans 600 0 0 0 serial_clock
port 34 nsew
flabel metal3 s 14000 13472 34000 13592 0 FreeSans 600 0 0 0 serial_clock_out
port 35 nsew
flabel metal3 s 14000 13880 34000 14000 0 FreeSans 600 0 0 0 serial_data_in
port 36 nsew
flabel metal3 s 14000 14288 34000 14408 0 FreeSans 600 0 0 0 serial_data_out
port 37 nsew
flabel metal3 s 14000 14696 34000 14816 0 FreeSans 600 0 0 0 serial_load
port 38 nsew
flabel metal3 s 14000 15104 34000 15224 0 FreeSans 600 0 0 0 serial_load_out
port 39 nsew
flabel metal3 s 14000 15512 34000 15632 0 FreeSans 600 0 0 0 user_gpio_in
port 40 nsew
flabel metal3 s 14000 15920 34000 16040 0 FreeSans 600 0 0 0 user_gpio_oeb
port 41 nsew
flabel metal3 s 14000 16328 34000 16448 0 FreeSans 600 0 0 0 user_gpio_out
port 42 nsew
flabel metal4 s 2560 4893 2880 15824 0 FreeSans 2400 90 0 0 vccd
port 43 nsew
flabel metal4 s 7560 928 7880 15824 0 FreeSans 2400 90 0 0 vccd
port 43 nsew
flabel metal5 s 872 928 9892 1248 0 FreeSans 3200 0 0 0 vccd
port 43 nsew
flabel metal5 s 872 4928 9892 5248 0 FreeSans 3200 0 0 0 vccd
port 43 nsew
flabel metal5 s 872 8928 9892 9248 0 FreeSans 3200 0 0 0 vccd
port 43 nsew
flabel metal5 s 872 12928 9892 13248 0 FreeSans 3200 0 0 0 vccd
port 43 nsew
flabel metal4 s 4560 1040 4880 15824 0 FreeSans 2400 90 0 0 vccd1
port 44 nsew
flabel metal4 s 9560 1040 9880 15824 0 FreeSans 2400 90 0 0 vccd1
port 44 nsew
flabel metal5 s 872 2928 9892 3248 0 FreeSans 3200 0 0 0 vccd1
port 44 nsew
flabel metal5 s 872 6928 9892 7248 0 FreeSans 3200 0 0 0 vccd1
port 44 nsew
flabel metal5 s 872 10928 9892 11248 0 FreeSans 3200 0 0 0 vccd1
port 44 nsew
flabel metal5 s 872 14928 9892 15248 0 FreeSans 3200 0 0 0 vccd1
port 44 nsew
flabel metal4 s 3560 1040 3880 15824 0 FreeSans 2400 90 0 0 vssd
port 45 nsew
flabel metal4 s 8560 1040 8880 15824 0 FreeSans 2400 90 0 0 vssd
port 45 nsew
flabel metal5 s 872 1928 9892 2248 0 FreeSans 3200 0 0 0 vssd
port 45 nsew
flabel metal5 s 872 5928 9892 6248 0 FreeSans 3200 0 0 0 vssd
port 45 nsew
flabel metal5 s 872 9928 9892 10248 0 FreeSans 3200 0 0 0 vssd
port 45 nsew
flabel metal5 s 872 13928 9892 14248 0 FreeSans 3200 0 0 0 vssd
port 45 nsew
flabel metal4 s 5560 1040 5880 15824 0 FreeSans 2400 90 0 0 vssd1
port 46 nsew
flabel metal5 s 872 3928 9892 4248 0 FreeSans 3200 0 0 0 vssd1
port 46 nsew
flabel metal3 s 14000 4496 34000 4616 0 FreeSans 600 0 0 0 zero
port 47 nsew
<< properties >>
string FIXED_BBOX 0 0 34000 17000
<< end >>
